////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/// TSMC Library/IP Product
/// Filename: tcbn28hpcplusbwp7t30p140hvt.v
/// Technology: CLN28HT
/// Product Type: Standard Cell
/// Product Name: tcbn28hpcplusbwp7t30p140hvt
/// Version: 110a
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////
///  STATEMENT OF USE
///
///  This information contains confidential and proprietary information of TSMC.
///  No part of this information may be reproduced, transmitted, transcribed,
///  stored in a retrieval system, or translated into any human or computer
///  language, in any form or by any means, electronic, mechanical, magnetic,
///  optical, chemical, manual, or otherwise, without the prior written permission
///  of TSMC.  This information was prepared for informational purpose and is for
///  use by TSMC's customers only.  TSMC reserves the right to make changes in the
///  information at any time and without notice.
///
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps
`celldefine
module AN2D0BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2D8BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2OPTPAD12BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2OPTPAD1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2OPTPAD2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2OPTPAD4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN2OPTPAD8BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D0BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D1BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D2BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D4BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN3D8BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    and (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D0BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D1BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D2BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D4BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AN4D8BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    and (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ANTENNABWP7T30P140HVT (I);
    input I;
    buf (I_buf, I);

endmodule
`endcelldefine

`celldefine
module AO211D0BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D1BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D2BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO211D4BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D0BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D1BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D2BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO21D4BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    and (I0_out, A1, A2);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D0BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D1BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D2BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO221D4BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D0BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D1BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D2BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO222D4BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    and (I2_out, C1, C2);
    or (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D0BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D1BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D2BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO22D4BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D0BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D1BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D2BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO31D4BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    and (I0_out, A1, A2, A3);
    or (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D0BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D1BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D2BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO32D4BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D0BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D1BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D2BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AO33D4BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    and (I0_out, A1, A2, A3);
    and (I1_out, B1, B2, B3);
    or (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D0BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D1BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D2BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211D4BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211OPTBD12BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211OPTBD1BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211OPTBD2BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211OPTBD4BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211OPTBD6BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI211OPTBD8BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    and (I0_out, A1, A2);
    or (I2_out, I0_out, B, C);
    not (ZN, I2_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D0BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21D4BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21OPTBD12BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21OPTBD1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21OPTBD2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21OPTBD4BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21OPTBD6BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI21OPTBD8BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D0BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D1BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D2BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI221D4BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D0BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D1BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D2BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI222D4BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, C1, C2);
    and (I2_out, B1, B2);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C2 == 1'b1)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && C1 == 1'b1)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D0BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22D4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22OPTPBD12BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22OPTPBD1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22OPTPBD2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22OPTPBD4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22OPTPBD6BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI22OPTPBD8BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D0BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D1BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D2BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI31D4BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    and (I0_out, A1, A2, A3);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D0BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D1BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D2BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI32D4BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    and (I0_out, B1, B2);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D0BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D1BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D2BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module AOI33D4BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    and (I0_out, B1, B2, B3);
    and (I1_out, A1, A2, A3);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B3 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BHDBWP7T30P140HVT (Z);
    inout Z;
    not (weak0, weak1) (Z, Z_buf);
    not                (Z_buf, Z);

endmodule
`endcelldefine

`celldefine
module BOUNDARY_LEFTBWP7T30P140;
    // No function
endmodule
`endcelldefine

`celldefine
module BOUNDARY_RIGHTBWP7T30P140;
    // No function
endmodule
`endcelldefine

`celldefine
module BUFFD0BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD12BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD16BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD20BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD3BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD6BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFFD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD12BWP7T30P140HVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD16BWP7T30P140HVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD4BWP7T30P140HVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD6BWP7T30P140HVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module BUFTD8BWP7T30P140HVT (I, OE, Z);
    input I, OE;
    output Z;
    bufif1 (Z, I, OE);

  specify
    (I => Z) = (0, 0);
    (OE => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D0BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKAN2D8BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD0BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD12BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD16BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD20BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD3BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD6BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKBD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKLHQD12BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD16BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD1BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD2BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD3BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD4BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD6BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLHQD8BWP7T30P140HVT ( Q, TE, CPN, E );
    input TE, CPN, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, CPN_d, E_d;
        buf (_TE, TE_d);
        buf (_CPN, CPN_d);
        buf (_E, E_d);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `else 
        buf (_TE, TE);
        buf (_CPN, CPN);
        buf (_E, E);
        or (_G001, _E, _TE);
        tsmc_dla (_enl, _G001, _CPN, 1'b1, 1'b1, notifier);
        not (_enlb, _enl);
        or (Q, _enlb, _CPN);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b0 && TE == 1'b0)
    (posedge CPN => (Q+:1'b1)) = (0, 0);
    if (E == 1'b1 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CPN => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CPN => Q) = (0, 0);
    $width (posedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CPN_d, E_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CPN_d, TE_d);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CPN_d, TE_d);
  `else
    $setuphold (negedge CPN &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD12BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD16BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD1BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD20BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD2BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD3BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD4BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD6BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQD8BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQOPTMAD12BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQOPTMAD4BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKLNQOPTMAD8BWP7T30P140HVT (TE, E, CP, Q);
    input TE, E, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire TE_d, E_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        or (D_i, E_d, TE_d);
        not (CPB, CP_d);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP_d);
    `else 
        pullup (CDN);
        pullup (SDN);
        or (D_i, E, TE);
        not (CPB, CP);
        tsmc_dla (Q_buf, D_i, CPB, CDN, SDN, notifier);
        and (Q, Q_buf, CP);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (nTE_SDFCHK, nTE, 1'b1);
    tsmc_xbuf (nE_SDFCHK, nE, 1'b1);
    tsmc_xbuf (E_TE_SDFCHK, E_TE, 1'b1);
    tsmc_xbuf (E_nTE_SDFCHK, E_nTE, 1'b1);
    tsmc_xbuf (nE_TE_SDFCHK, nE_TE, 1'b1);
    tsmc_xbuf (nE_nTE_SDFCHK, nE_nTE, 1'b1);
    not (nTE, TE);
    not (nE, E);
    and (E_TE, E, TE);
    and (E_nTE, E, nTE);
    and (nE_TE, nE, TE);
    and (nE_nTE, nE, nTE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (E_int_not, E_d);
      not  (TE_int_not, TE_d);
    `else
      not  (E_int_not, E);
      not  (TE_int_not, TE);
    `endif
    buf  (E_check, TE_int_not);
    buf  (TE_check, E_int_not);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);
    tsmc_xbuf (TE_DEFCHK, TE_check, 1'b1);

  specify
    if (E == 1'b1 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b1 && TE == 1'b0)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b1)
    (CP => Q) = (0, 0);
    if (E == 1'b0 && TE == 1'b0)
    (negedge CP => (Q+:1'b0)) = (0, 0);
    $width (posedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_TE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& E_nTE_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_TE_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nE_nTE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier,,, CP_d, E_d);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier,,, CP_d, TE_d);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier,,, CP_d, TE_d);
  `else
    $setuphold (posedge CP &&& nTE_SDFCHK, posedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nTE_SDFCHK, negedge E , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, posedge TE , 0, 0, notifier);
    $setuphold (posedge CP &&& nE_SDFCHK, negedge TE , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module CKMUX2D0BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D1BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D2BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKMUX2D4BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND0BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND12BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND16BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND1BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND20BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D0BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D3BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND2D8BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND3BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND4BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND6BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKND8BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D0BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module CKXOR2D4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCAP16BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP32BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP4BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP64BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCAP8BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module DCCKBD12BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKBD16BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKBD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKBD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKND12BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKND16BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKND20BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKND4BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DCCKND8BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL025D1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL050MD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL075MD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL100MD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL150MD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL200MD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DEL250MD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module DFCND1BWP7T30P140HVT (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCND2BWP7T30P140HVT (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCND4BWP7T30P140HVT (D, CP, CDN, Q, QN);
    input D, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD1BWP7T30P140HVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD2BWP7T30P140HVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCNQD4BWP7T30P140HVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND1BWP7T30P140HVT (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CP_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND2BWP7T30P140HVT (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CP_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSND4BWP7T30P140HVT (D, CP, CDN, SDN, Q, QN);
    input D, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CP_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD1BWP7T30P140HVT (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CP_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD2BWP7T30P140HVT (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CP_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFCSNQD4BWP7T30P140HVT (D, CP, CDN, SDN, Q);
    input D, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SDFCHK, CP_D_SDN, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SDFCHK, CP_nD_SDN, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SDFCHK, nCP_D_SDN, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SDFCHK, nCP_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CP_D_SDFCHK, CDN_CP_D, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SDFCHK, CDN_CP_nD, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SDFCHK, CDN_nCP_D, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SDFCHK, CDN_nCP_nD, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D_SDN, CP, D, SDN);
    and (CP_nD_SDN, CP, nD, SDN);
    and (nCP_D_SDN, nCP, D, SDN);
    and (nCP_nD_SDN, nCP, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CP_D, CDN, CP, D);
    and (CDN_CP_nD, CDN, CP, nD);
    and (CDN_nCP_D, CDN, nCP, D);
    and (CDN_nCP_nD, CDN, nCP, nD);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CP_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge CP &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge CP &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD1BWP7T30P140HVT (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD2BWP7T30P140HVT (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFD4BWP7T30P140HVT (D, CP, Q, QN);
    input D, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND1BWP7T30P140HVT (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, CN_d);
    `else
      buf  (D_check, CN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND2BWP7T30P140HVT (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, CN_d);
    `else
      buf  (D_check, CN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCND4BWP7T30P140HVT (D, CP, CN, Q, QN);
    input D, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, CN_d);
    `else
      buf  (D_check, CN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    (posedge CP => (QN-:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD1BWP7T30P140HVT (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, CN_d);
    `else
      buf  (D_check, CN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD2BWP7T30P140HVT (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, CN_d);
    `else
      buf  (D_check, CN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCNQD4BWP7T30P140HVT (D, CP, CN, Q);
    input D, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN_d, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D_i, CN, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CN_SDFCHK, CN, 1'b1);
    tsmc_xbuf (CN_D_SDFCHK, CN_D, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    tsmc_xbuf (nCN_D_SDFCHK, nCN_D, 1'b1);
    tsmc_xbuf (nCN_nD_SDFCHK, nCN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    and (CN_D, CN, D);
    and (CN_nD, CN, nD);
    and (nCN_D, nCN, D);
    and (nCN_nD, nCN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, CN_d);
    `else
      buf  (D_check, CN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D)))) = (0, 0);
    $width (posedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SDFCHK, negedge D , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND1BWP7T30P140HVT (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D_i, CN_d, DS);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D_i, CN, DS);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SN_SDFCHK, CN_D_SN, 1'b1);
    tsmc_xbuf (CN_D_nSN_SDFCHK, CN_D_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSN_SDFCHK, CN_nD_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SN_SDFCHK, CN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_D_SN_SDFCHK, nCN_D_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSN_SDFCHK, nCN_D_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SN_SDFCHK, nCN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSN_SDFCHK, nCN_nD_nSN, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (CN_SN_SDFCHK, CN_SN, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SN, CN, D, SN);
    and (CN_D_nSN, CN, D, nSN);
    and (CN_nD_nSN, CN, nD, nSN);
    and (CN_nD_SN, CN, nD, SN);
    and (nCN_D_SN, nCN, D, SN);
    and (nCN_D_nSN, nCN, D, nSN);
    and (nCN_nD_SN, nCN, nD, SN);
    and (nCN_nD_nSN, nCN, nD, nSN);
    and (D_SN, D, SN);
    and (nD_nSN, nD, nSN);
    and (D_nSN, D, nSN);
    and (CN_SN, CN, SN);
    and (CN_nD, CN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (SN_check, CN_d);
      and  (D_check, SN_d, CN_d);
    `else
      buf  (SN_check, CN);
      and  (D_check, SN, CN);
    `endif
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND2BWP7T30P140HVT (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D_i, CN_d, DS);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D_i, CN, DS);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SN_SDFCHK, CN_D_SN, 1'b1);
    tsmc_xbuf (CN_D_nSN_SDFCHK, CN_D_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSN_SDFCHK, CN_nD_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SN_SDFCHK, CN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_D_SN_SDFCHK, nCN_D_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSN_SDFCHK, nCN_D_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SN_SDFCHK, nCN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSN_SDFCHK, nCN_nD_nSN, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (CN_SN_SDFCHK, CN_SN, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SN, CN, D, SN);
    and (CN_D_nSN, CN, D, nSN);
    and (CN_nD_nSN, CN, nD, nSN);
    and (CN_nD_SN, CN, nD, SN);
    and (nCN_D_SN, nCN, D, SN);
    and (nCN_D_nSN, nCN, D, nSN);
    and (nCN_nD_SN, nCN, nD, SN);
    and (nCN_nD_nSN, nCN, nD, nSN);
    and (D_SN, D, SN);
    and (nD_nSN, nD, nSN);
    and (D_nSN, D, nSN);
    and (CN_SN, CN, SN);
    and (CN_nD, CN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (SN_check, CN_d);
      and  (D_check, SN_d, CN_d);
    `else
      buf  (SN_check, CN);
      and  (D_check, SN, CN);
    `endif
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKCSND4BWP7T30P140HVT (D, CP, CN, SN, Q, QN);
    input D, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D_i, CN_d, DS);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D_i, CN, DS);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SN_SDFCHK, CN_D_SN, 1'b1);
    tsmc_xbuf (CN_D_nSN_SDFCHK, CN_D_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSN_SDFCHK, CN_nD_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SN_SDFCHK, CN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_D_SN_SDFCHK, nCN_D_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSN_SDFCHK, nCN_D_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SN_SDFCHK, nCN_nD_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSN_SDFCHK, nCN_nD_nSN, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (CN_SN_SDFCHK, CN_SN, 1'b1);
    tsmc_xbuf (CN_nD_SDFCHK, CN_nD, 1'b1);
    not (nD, D);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SN, CN, D, SN);
    and (CN_D_nSN, CN, D, nSN);
    and (CN_nD_nSN, CN, nD, nSN);
    and (CN_nD_SN, CN, nD, SN);
    and (nCN_D_SN, nCN, D, SN);
    and (nCN_D_nSN, nCN, D, nSN);
    and (nCN_nD_SN, nCN, nD, SN);
    and (nCN_nD_nSN, nCN, nD, nSN);
    and (D_SN, D, SN);
    and (nD_nSN, nD, nSN);
    and (D_nSN, D, nSN);
    and (CN_SN, CN, SN);
    and (CN_nD, CN, nD);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (SN_check, CN_d);
      and  (D_check, SN_d, CN_d);
    `else
      buf  (SN_check, CN);
      and  (D_check, SN, CN);
    `endif
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((CN && D) || (CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND1BWP7T30P140HVT (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D_i, S, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D_i, S, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_SDFCHK, SN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (nD_SN_SDFCHK, nD_SN, 1'b1);
    not (nD, D);
    not (nSN, SN);
    and (D_SN, D, SN);
    and (D_nSN, D, nSN);
    and (nD_nSN, nD, nSN);
    and (nD_SN, nD, SN);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, SN_d);
    `else
      buf  (D_check, SN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND2BWP7T30P140HVT (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D_i, S, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D_i, S, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_SDFCHK, SN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (nD_SN_SDFCHK, nD_SN, 1'b1);
    not (nD, D);
    not (nSN, SN);
    and (D_SN, D, SN);
    and (D_nSN, D, nSN);
    and (nD_nSN, nD, nSN);
    and (nD_SN, nD, SN);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, SN_d);
    `else
      buf  (D_check, SN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFKSND4BWP7T30P140HVT (D, CP, SN, Q, QN);
    input D, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D_i, S, D_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D_i, S, D);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SN_SDFCHK, SN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SN_SDFCHK, D_SN, 1'b1);
    tsmc_xbuf (D_nSN_SDFCHK, D_nSN, 1'b1);
    tsmc_xbuf (nD_nSN_SDFCHK, nD_nSN, 1'b1);
    tsmc_xbuf (nD_SN_SDFCHK, nD_SN, 1'b1);
    not (nD, D);
    not (nSN, SN);
    and (D_SN, D, SN);
    and (D_nSN, D, nSN);
    and (nD_nSN, nD, nSN);
    and (nD_SN, nD, SN);


  // Timing logics defined for default constraint check
    `ifdef NTC
      buf  (D_check, SN_d);
    `else
      buf  (D_check, SN);
    `endif
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((D) || (!(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((D) || (!(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFMD1BWP7T30P140HVT (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      buf  (DA_check, SA_d);
    `else
      not  (SA_int_not, SA);
      buf  (DA_check, SA);
    `endif
    buf  (DB_check, SA_int_not);
    pullup  (CP_check);
    pullup  (SA_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);

  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFMD2BWP7T30P140HVT (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      buf  (DA_check, SA_d);
    `else
      not  (SA_int_not, SA);
      buf  (DA_check, SA);
    `endif
    buf  (DB_check, SA_int_not);
    pullup  (CP_check);
    pullup  (SA_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);

  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFMD4BWP7T30P140HVT (DA, DB, SA, CP, Q, QN);
    input DA, DB, SA, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      buf  (DA_check, SA_d);
    `else
      not  (SA_int_not, SA);
      buf  (DA_check, SA);
    `endif
    buf  (DB_check, SA_int_not);
    pullup  (CP_check);
    pullup  (SA_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);

  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    (posedge CP => (QN-:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFMQD1BWP7T30P140HVT (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      buf  (DA_check, SA_d);
    `else
      not  (SA_int_not, SA);
      buf  (DA_check, SA);
    `endif
    buf  (DB_check, SA_int_not);
    pullup  (CP_check);
    pullup  (SA_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);

  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFMQD2BWP7T30P140HVT (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      buf  (DA_check, SA_d);
    `else
      not  (SA_int_not, SA);
      buf  (DA_check, SA);
    `endif
    buf  (DB_check, SA_int_not);
    pullup  (CP_check);
    pullup  (SA_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);

  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFMQD4BWP7T30P140HVT (DA, DB, SA, CP, Q);
    input DA, DB, SA, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_dff (Q_buf, D, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SDFCHK, DA_DB_SA, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SDFCHK, DA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SDFCHK, DA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SDFCHK, nDA_DB_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SDFCHK, DA_nDB_nSA, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SDFCHK, nDA_DB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SDFCHK, nDA_nDB_SA, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SDFCHK, nDA_nDB_nSA, 1'b1);
    tsmc_xbuf (DB_SA_SDFCHK, DB_SA, 1'b1);
    tsmc_xbuf (nDB_SA_SDFCHK, nDB_SA, 1'b1);
    tsmc_xbuf (DA_nSA_SDFCHK, DA_nSA, 1'b1);
    tsmc_xbuf (nDA_nSA_SDFCHK, nDA_nSA, 1'b1);
    tsmc_xbuf (DA_nDB_SDFCHK, DA_nDB, 1'b1);
    tsmc_xbuf (nDA_DB_SDFCHK, nDA_DB, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    and (DA_DB_SA, DA, DB, SA);
    and (DA_DB_nSA, DA, DB, nSA);
    and (DA_nDB_SA, DA, nDB, SA);
    and (nDA_DB_nSA, nDA, DB, nSA);
    and (DA_nDB_nSA, DA, nDB, nSA);
    and (nDA_DB_SA, nDA, DB, SA);
    and (nDA_nDB_SA, nDA, nDB, SA);
    and (nDA_nDB_nSA, nDA, nDB, nSA);
    and (DB_SA, DB, SA);
    and (nDB_SA, nDB, SA);
    and (DA_nSA, DA, nSA);
    and (nDA_nSA, nDA, nSA);
    and (DA_nDB, DA, nDB);
    and (nDA_DB, nDA, DB);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      buf  (DA_check, SA_d);
    `else
      not  (SA_int_not, SA);
      buf  (DA_check, SA);
    `endif
    buf  (DB_check, SA_int_not);
    pullup  (CP_check);
    pullup  (SA_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);

  specify
    (posedge CP => (Q+:((DA && DB) || (DA && !(DB) && SA) || (!(DA) && DB && !(SA))))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
  `else
    $setuphold (posedge CP &&& DB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SDFCHK, negedge SA , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND1BWP7T30P140HVT (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CPN_d;
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CPN_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND2BWP7T30P140HVT (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CPN_d;
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CPN_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCND4BWP7T30P140HVT (D, CPN, CDN, Q, QN);
    input D, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CPN_d;
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CPN_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge CPN &&& D_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND1BWP7T30P140HVT (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SDFCHK, CPN_D_SDN, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SDFCHK, CPN_nD_SDN, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SDFCHK, nCPN_D_SDN, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SDFCHK, nCPN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SDFCHK, CDN_CPN_D, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SDFCHK, CDN_CPN_nD, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SDFCHK, CDN_nCPN_D, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SDFCHK, CDN_nCPN_nD, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D_SDN, CPN, D, SDN);
    and (CPN_nD_SDN, CPN, nD, SDN);
    and (nCPN_D_SDN, nCPN, D, SDN);
    and (nCPN_nD_SDN, nCPN, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CPN_D, CDN, CPN, D);
    and (CDN_CPN_nD, CDN, CPN, nD);
    and (CDN_nCPN_D, CDN, nCPN, D);
    and (CDN_nCPN_nD, CDN, nCPN, nD);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CPN_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND2BWP7T30P140HVT (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SDFCHK, CPN_D_SDN, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SDFCHK, CPN_nD_SDN, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SDFCHK, nCPN_D_SDN, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SDFCHK, nCPN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SDFCHK, CDN_CPN_D, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SDFCHK, CDN_CPN_nD, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SDFCHK, CDN_nCPN_D, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SDFCHK, CDN_nCPN_nD, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D_SDN, CPN, D, SDN);
    and (CPN_nD_SDN, CPN, nD, SDN);
    and (nCPN_D_SDN, nCPN, D, SDN);
    and (nCPN_nD_SDN, nCPN, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CPN_D, CDN, CPN, D);
    and (CDN_CPN_nD, CDN, CPN, nD);
    and (CDN_nCPN_D, CDN, nCPN, D);
    and (CDN_nCPN_nD, CDN, nCPN, nD);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CPN_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNCSND4BWP7T30P140HVT (D, CPN, CDN, SDN, Q, QN);
    input D, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SDFCHK, CPN_D_SDN, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SDFCHK, CPN_nD_SDN, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SDFCHK, nCPN_D_SDN, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SDFCHK, nCPN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SDFCHK, CDN_CPN_D, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SDFCHK, CDN_CPN_nD, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SDFCHK, CDN_nCPN_D, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SDFCHK, CDN_nCPN_nD, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (CPN_D_SDN, CPN, D, SDN);
    and (CPN_nD_SDN, CPN, nD, SDN);
    and (nCPN_D_SDN, nCPN, D, SDN);
    and (nCPN_nD_SDN, nCPN, nD, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_CPN_D, CDN, CPN, D);
    and (CDN_CPN_nD, CDN, CPN, nD);
    and (CDN_nCPN_D, CDN, nCPN, D);
    and (CDN_nCPN_nD, CDN, nCPN, nD);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (CPN_check, CDN_i, SDN_i);
    and  (D_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge CPN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge CPN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND1BWP7T30P140HVT (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CPN_check);
    pullup  (D_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND2BWP7T30P140HVT (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CPN_check);
    pullup  (D_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFND4BWP7T30P140HVT (D, CPN, Q, QN);
    input D, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CPN_check);
    pullup  (D_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    $width (posedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CPN_d, D_d);
  `else
    $setuphold (negedge CPN &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (negedge CPN &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND1BWP7T30P140HVT (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        pullup (CDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);


  // Timing logics defined for default constraint check
    buf  (CPN_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND2BWP7T30P140HVT (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        pullup (CDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);


  // Timing logics defined for default constraint check
    buf  (CPN_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFNSND4BWP7T30P140HVT (D, CPN, SDN, Q, QN);
    input D, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CPN_d;
        pullup (CDN);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_d, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (CP, CPN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CPN_D_SDFCHK, CPN_D, 1'b1);
    tsmc_xbuf (CPN_nD_SDFCHK, CPN_nD, 1'b1);
    tsmc_xbuf (nCPN_D_SDFCHK, nCPN_D, 1'b1);
    tsmc_xbuf (nCPN_nD_SDFCHK, nCPN_nD, 1'b1);
    not (nD, D);
    not (nCPN, CPN);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CPN_D, CPN, D);
    and (CPN_nD, CPN, nD);
    and (nCPN_D, nCPN, D);
    and (nCPN_nD, nCPN, nD);


  // Timing logics defined for default constraint check
    buf  (CPN_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (negedge CPN => (Q+:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:D)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge CPN &&& nD_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD1BWP7T30P140HVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD2BWP7T30P140HVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFQD4BWP7T30P140HVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND1BWP7T30P140HVT (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND2BWP7T30P140HVT (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSND4BWP7T30P140HVT (D, CP, SDN, Q, QN);
    input D, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD1BWP7T30P140HVT (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD2BWP7T30P140HVT (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module DFSNQD4BWP7T30P140HVT (D, CP, SDN, Q);
    input D, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, CP_d;
        pullup (CDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, SDN_i);
    buf  (D_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
      $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge CP &&& nD_SDFCHK, 0, notifier);
    $hold (posedge CP &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module FA1D0BWP7T30P140HVT (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D1BWP7T30P140HVT (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D2BWP7T30P140HVT (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1D4BWP7T30P140HVT (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1OPTCD1BWP7T30P140HVT (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FA1OPTSD1BWP7T30P140HVT (A, B, CI, S, CO);
    input A, B, CI;
    output S, CO;
    xor (I0_out, A, B);
    xor (S, I0_out, CI);
    and (I1_out, A, B);
    and (I2_out, B, CI);
    and (I3_out, A, CI);
    or (CO, I1_out, I2_out, I3_out);

  specify
    if (B == 1'b1 && CI == 1'b0)
    (A => CO) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => CO) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => CO) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => CO) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => CO) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => CO) = (0, 0);
    if (B == 1'b1 && CI == 1'b1)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1 && CI == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b0 && CI == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1 && CI == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b0 && CI == 1'b1)
    (B => S) = (0, 0);
    if (A == 1'b1 && B == 1'b1)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (CI => S) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (CI => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module FILL16BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module FILL2BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module FILL32BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module FILL3BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module FILL4BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module FILL64BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module FILL8BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GAN2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2MCOD1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAN2MCOD2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    and (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI21D1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI21D2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI21MCOD1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI21MCOD2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    and (I0_out, A1, A2);
    or (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI22D1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GAOI22MCOD1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    and (I1_out, B1, B2);
    or (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD3BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFMCOD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFMCOD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFMCOD3BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFMCOD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GBUFFMCOD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GDCAP10BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP10MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP12BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP12MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP2BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP2MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP3BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP3MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP4BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAP4MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAPBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDCAPMCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GDFCNQD1BWP7T30P140HVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GDFCNQMCOD1BWP7T30P140HVT (D, CP, CDN, Q);
    input D, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, CP_d;
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (CP_D_SDFCHK, CP_D, 1'b1);
    tsmc_xbuf (CP_nD_SDFCHK, CP_nD, 1'b1);
    tsmc_xbuf (nCP_D_SDFCHK, nCP_D, 1'b1);
    tsmc_xbuf (nCP_nD_SDFCHK, nCP_nD, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nCP, CP);
    and (CP_D, CP, D);
    and (CP_nD, CP, nD);
    and (nCP_D, nCP, D);
    and (nCP_nD, nCP, nD);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (CP_check, CDN_i);
    buf  (D_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge CP &&& D_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GDFQD1BWP7T30P140HVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GDFQMCOD1BWP7T30P140HVT (D, CP, Q);
    input D, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D_d, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dff (Q_buf, D, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  // Timing logics defined for default constraint check
    pullup  (CP_check);
    pullup  (D_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:D)) = (0, 0);
    $width (posedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier,,, CP_d, D_d);
  `else
    $setuphold (posedge CP &&& D_DEFCHK, posedge D, 0, 0, notifier);
    $setuphold (posedge CP &&& D_DEFCHK, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GFILL10BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL10MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL12BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL12MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL2BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL2MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL3BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL3MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL4BWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILL4MCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILLBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GFILLMCOBWP7T30P140HVT;
    // No function
endmodule
`endcelldefine

`celldefine
module GINVD1BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD2BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD3BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD4BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVD8BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVMCOD1BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVMCOD2BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVMCOD3BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVMCOD4BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GINVMCOD8BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2D1BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2D2BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2MCOD1BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2MCOD2BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2ND1BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2ND2BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2NMCOD1BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GMUX2NMCOD2BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D3BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2D4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2MCOD1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2MCOD2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2MCOD3BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND2MCOD4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3D1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3D2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3MCOD1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GND3MCOD2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2MCOD1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR2MCOD2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR3D1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR3D2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR3MCOD1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GNR3MCOD2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOAI21D1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOAI21D2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOAI21MCOD1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOAI21MCOD2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2MCOD1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GOR2MCOD2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GSDFCNQD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GSDFCNQMCOD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module GTIEHBWP7T30P140HVT (Z);
    output Z;
    buf (Z, 1'b1);

endmodule
`endcelldefine

`celldefine
module GTIEHMCOBWP7T30P140HVT (Z);
    output Z;
    buf (Z, 1'b1);

endmodule
`endcelldefine

`celldefine
module GTIELBWP7T30P140HVT (ZN);
    output ZN;
    buf (ZN, 1'b0);

endmodule
`endcelldefine

`celldefine
module GTIELMCOBWP7T30P140HVT (ZN);
    output ZN;
    buf (ZN, 1'b0);

endmodule
`endcelldefine

`celldefine
module GXNR2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXNR2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXNR2MCOD1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXNR2MCOD2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2MCOD1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module GXOR2MCOD2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D0BWP7T30P140HVT (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D1BWP7T30P140HVT (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D2BWP7T30P140HVT (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module HA1D4BWP7T30P140HVT (A, B, S, CO);
    input A, B;
    output S, CO;
    xor (S, A, B);
    and (CO, A, B);

  specify
    (A => CO) = (0, 0);
    (B => CO) = (0, 0);
    if (B == 1'b0)
    (A => S) = (0, 0);
    if (B == 1'b1)
    (A => S) = (0, 0);
    if (A == 1'b0)
    (B => S) = (0, 0);
    if (A == 1'b1)
    (B => S) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D0BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D1BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D2BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2D4BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2OPTPAD12BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2OPTPAD1BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2OPTPAD2BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2OPTPAD4BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND2OPTPAD8BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D0BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D1BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D2BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND3D4BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D0BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D1BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D2BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module IND4D4BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    and (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D0BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D1BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D2BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2D4BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2OPTPAD12BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2OPTPAD1BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2OPTPAD2BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2OPTPAD4BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR2OPTPAD8BWP7T30P140HVT (A1, B1, ZN);
    input A1, B1;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D0BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D1BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D2BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR3D4BWP7T30P140HVT (A1, B1, B2, ZN);
    input A1, B1, B2;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D0BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D1BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D2BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INR4D4BWP7T30P140HVT (A1, B1, B2, B3, ZN);
    input A1, B1, B2, B3;
    output ZN;
    not (I0_out, A1);
    or (I1_out, I0_out, B1, B2, B3);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (B1 => ZN) = (0, 0);
    (B2 => ZN) = (0, 0);
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD0BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD12BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD16BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD1BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD20BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD2BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD3BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD4BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD6BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module INVD8BWP7T30P140HVT (I, ZN);
    input I;
    output ZN;
    not (ZN, I);

  specify
    (I => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LHCND1BWP7T30P140HVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCND2BWP7T30P140HVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCND4BWP7T30P140HVT (D, E, CDN, Q, QN);
    input D, E, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD1BWP7T30P140HVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD2BWP7T30P140HVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCNQD4BWP7T30P140HVT (D, E, CDN, Q);
    input D, E, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, E_d;
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
    `else
      $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, negedge E &&& D_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND1BWP7T30P140HVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND2BWP7T30P140HVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSND4BWP7T30P140HVT (D, E, CDN, SDN, Q, QN);
    input D, E, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD1BWP7T30P140HVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => Q) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD2BWP7T30P140HVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => Q) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHCSNQD4BWP7T30P140HVT (D, E, CDN, SDN, Q);
    input D, E, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        tsmc_dla (Q_buf, D_d, E_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_nE_SDN_SDFCHK, D_nE_SDN, 1'b1);
    tsmc_xbuf (nD_nE_SDN_SDFCHK, nD_nE_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_nE_SDFCHK, CDN_D_nE, 1'b1);
    tsmc_xbuf (CDN_nD_nE_SDFCHK, CDN_nD_nE, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_nE_SDN, D, nE, SDN);
    and (nD_nE_SDN, nD, nE, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_nE, CDN, D, nE);
    and (CDN_nD_nE, CDN, nD, nE);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    if (D == 1'b1 && E == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && E == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && E == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && E == 1'b0)
    (SDN => Q) = (0, 0);
    $width (negedge CDN &&& D_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_nE_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, E_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
      $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_nE_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_nE_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, negedge E &&& D_SDN_SDFCHK, 0, notifier);
    $hold (negedge E &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, negedge E &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD1BWP7T30P140HVT (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD2BWP7T30P140HVT (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHD4BWP7T30P140HVT (D, E, Q, QN);
    input D, E;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHQD1BWP7T30P140HVT (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHQD2BWP7T30P140HVT (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHQD4BWP7T30P140HVT (D, E, Q);
    input D, E;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, E_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    $width (posedge E &&& D_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge E, posedge D, 0, 0, notifier,,, E_d, D_d);
    $setuphold (negedge E, negedge D, 0, 0, notifier,,, E_d, D_d);
  `else
    $setuphold (negedge E, posedge D, 0, 0, notifier);
    $setuphold (negedge E, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND1BWP7T30P140HVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    ifnone (posedge SDN => (QN+:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND2BWP7T30P140HVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    ifnone (posedge SDN => (QN+:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSND4BWP7T30P140HVT (D, E, SDN, Q, QN);
    input D, E, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (posedge E => (QN-:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    ifnone (posedge SDN => (QN+:1'b1)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD1BWP7T30P140HVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD2BWP7T30P140HVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LHSNQD4BWP7T30P140HVT (D, E, SDN, Q);
    input D, E, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, E_d;
        pullup (CDN);
        tsmc_dla (Q_buf, D_d, E_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_nE_SDFCHK, D_nE, 1'b1);
    tsmc_xbuf (nD_nE_SDFCHK, nD_nE, 1'b1);
    not (nD, D);
    not (nE, E);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_nE, D, nE);
    and (nD_nE, nD, nE);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (E_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (E_DEFCHK, E_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (posedge E => (Q+:D)) = (0, 0);
    if (D == 1'b1 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && E == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    $width (posedge E &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (posedge E &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_nE_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_nE_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, E_d);
    `else
      $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, E_d, D_d);
      $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, E_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
      $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge E &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge E &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, negedge E &&& nD_SDFCHK, 0, notifier);
    $hold (negedge E &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND1BWP7T30P140HVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND2BWP7T30P140HVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCND4BWP7T30P140HVT (D, EN, CDN, Q, QN);
    input D, EN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD1BWP7T30P140HVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD2BWP7T30P140HVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCNQD4BWP7T30P140HVT (D, EN, CDN, Q);
    input D, EN, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire D_d, EN_d;
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CDN_SDFCHK, CDN, 1'b1);
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_D_SDFCHK, CDN_D, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_D, CDN, D);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    buf  (D_check, CDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge CDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& CDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDFCHK, posedge EN &&& D_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND1BWP7T30P140HVT (D, EN, CDN, SDN, Q, QN);
    input D, EN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND2BWP7T30P140HVT (D, EN, CDN, SDN, Q, QN);
    input D, EN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSND4BWP7T30P140HVT (D, EN, CDN, SDN, Q, QN);
    input D, EN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    ifnone (posedge CDN => (QN-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD1BWP7T30P140HVT (D, EN, CDN, SDN, Q);
    input D, EN, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD2BWP7T30P140HVT (D, EN, CDN, SDN, Q);
    input D, EN, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNCSNQD4BWP7T30P140HVT (D, EN, CDN, SDN, Q);
    input D, EN, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (D_EN_SDN_SDFCHK, D_EN_SDN, 1'b1);
    tsmc_xbuf (nD_EN_SDN_SDFCHK, nD_EN_SDN, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SDFCHK, CDN_D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SDFCHK, CDN_nD_SDN, 1'b1);
    tsmc_xbuf (CDN_D_EN_SDFCHK, CDN_D_EN, 1'b1);
    tsmc_xbuf (CDN_nD_EN_SDFCHK, CDN_nD_EN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    tsmc_xbuf (CDN_SDN_SDFCHK, CDN_SDN, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (CDN_nD_SDFCHK, CDN_nD, 1'b1);
    not (nD, D);
    and (D_EN_SDN, D, EN, SDN);
    and (nD_EN_SDN, nD, EN, SDN);
    and (CDN_D_SDN, CDN, D, SDN);
    and (CDN_nD_SDN, CDN, nD, SDN);
    and (CDN_D_EN, CDN, D, EN);
    and (CDN_nD_EN, CDN, nD, EN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);
    and (CDN_SDN, CDN, SDN);
    and (D_SDN, D, SDN);
    and (CDN_nD, CDN, nD);


  // Timing logics defined for default constraint check
    and  (D_check, SDN_i, CDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    if (D == 1'b1 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b1 && EN == 1'b0 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1 && SDN == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    ifnone (posedge CDN => (Q+:1'b1)) = (0, 0);
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b1 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b1)
    (SDN => Q) = (0, 0);
    if (CDN == 1'b0 && D == 1'b0 && EN == 1'b0)
    (SDN => Q) = (0, 0);
    $width (negedge CDN &&& D_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nD_EN_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& CDN_nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recrem (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0,0, notifier, , , CDN_d, EN_d);
      $recrem (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
      $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& D_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nD_EN_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& CDN_SDN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& D_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nD_EN_SDFCHK, posedge SDN , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SDFCHK, posedge EN &&& D_SDN_SDFCHK, 0, notifier);
    $hold (posedge EN &&& D_SDN_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SDFCHK, posedge EN &&& CDN_nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& CDN_nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND1BWP7T30P140HVT (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND2BWP7T30P140HVT (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LND4BWP7T30P140HVT (D, EN, Q, QN);
    input D, EN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNQD1BWP7T30P140HVT (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNQD2BWP7T30P140HVT (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNQD4BWP7T30P140HVT (D, EN, Q);
    input D, EN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire D_d, EN_d;
        pullup (CDN);
        pullup (SDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDFCHK, D, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    not (nD, D);


  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    $width (negedge EN &&& D_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge EN, posedge D, 0, 0, notifier,,, EN_d, D_d);
    $setuphold (posedge EN, negedge D, 0, 0, notifier,,, EN_d, D_d);
  `else
    $setuphold (posedge EN, posedge D, 0, 0, notifier);
    $setuphold (posedge EN, negedge D, 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND1BWP7T30P140HVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    ifnone (posedge SDN => (QN+:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND2BWP7T30P140HVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    ifnone (posedge SDN => (QN+:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSND4BWP7T30P140HVT (D, EN, SDN, Q, QN);
    input D, EN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    (D => QN) = (0, 0);
    (negedge EN => (QN-:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    ifnone (posedge SDN => (QN+:1'b1)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD1BWP7T30P140HVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD2BWP7T30P140HVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module LNSNQD4BWP7T30P140HVT (D, EN, SDN, Q);
    input D, EN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire D_d, EN_d;
        pullup (CDN);
        not (E, EN_d);
        tsmc_dla (Q_buf, D_d, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        not (E, EN);
        tsmc_dla (Q_buf, D, E, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (SDN_SDFCHK, SDN, 1'b1);
    tsmc_xbuf (nD_SDFCHK, nD, 1'b1);
    tsmc_xbuf (D_SDN_SDFCHK, D_SDN, 1'b1);
    tsmc_xbuf (nD_SDN_SDFCHK, nD_SDN, 1'b1);
    tsmc_xbuf (D_EN_SDFCHK, D_EN, 1'b1);
    tsmc_xbuf (nD_EN_SDFCHK, nD_EN, 1'b1);
    not (nD, D);
    and (D_SDN, D, SDN);
    and (nD_SDN, nD, SDN);
    and (D_EN, D, EN);
    and (nD_EN, nD, EN);


  // Timing logics defined for default constraint check
    buf  (D_check, SDN_i);
    buf  (EN_check, SDN_i);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (EN_DEFCHK, EN_check, 1'b1);

  specify
    (D => Q) = (0, 0);
    (negedge EN => (Q+:D)) = (0, 0);
    if (D == 1'b1 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (D == 1'b0 && EN == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    ifnone (posedge SDN => (Q-:1'b0)) = (0, 0);
    $width (negedge EN &&& D_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge EN &&& nD_SDN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& D_EN_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nD_EN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recrem (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0,0, notifier, , , SDN_d, EN_d);
    `else
      $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier,,, EN_d, D_d);
      $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier,,, EN_d, D_d);
      $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
      $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge EN &&& SDN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge EN &&& SDN_SDFCHK, negedge D , 0, 0, notifier);
    $recovery (posedge SDN &&& nD_SDFCHK, posedge EN &&& nD_SDFCHK, 0, notifier);
    $hold (posedge EN &&& nD_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module MAOI222D0BWP7T30P140HVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D1BWP7T30P140HVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D2BWP7T30P140HVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI222D4BWP7T30P140HVT (A, B, C, ZN);
    input A, B, C;
    output ZN;
    and (I0_out, A, B);
    and (I1_out, B, C);
    and (I2_out, A, C);
    or (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (B == 1'b1 && C == 1'b0)
    (A => ZN) = (0, 0);
    if (B == 1'b0 && C == 1'b1)
    (A => ZN) = (0, 0);
    if (A == 1'b1 && C == 1'b0)
    (B => ZN) = (0, 0);
    if (A == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A == 1'b1 && B == 1'b0)
    (C => ZN) = (0, 0);
    if (A == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D0BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22D4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22OPTBD2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MAOI22OPTBD4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    and (I0_out, A1, A2);
    not (I1_out, I0_out);
    or (I2_out, B1, B2);
    and (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D0BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22D4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22OPTBD2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MOAI22OPTBD4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    not (I1_out, I0_out);
    and (I2_out, B1, B2);
    or (ZN, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D0BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D1BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D2BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2D4BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND0BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND1BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND2BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2ND4BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2NOPTND1BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2NOPTND2BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2NOPTND4BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2NOPTND6BWP7T30P140HVT (I0, I1, S, ZN);
    input I0, I1, S;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S);
    not (ZN, I0_out);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2OPTD1BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2OPTD2BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2OPTD4BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX2OPTD6BWP7T30P140HVT (I0, I1, S, Z);
    input I0, I1, S;
    output Z;
    tsmc_mux (Z, I0, I1, S);

  specify
    if (I1 == 1'b1 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && S == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && S == 1'b1)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1)
    (S => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0)
    (S => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D0BWP7T30P140HVT (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D1BWP7T30P140HVT (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D2BWP7T30P140HVT (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3D4BWP7T30P140HVT (I0, I1, I2, S0, S1, Z);
    input I0, I1, I2, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (Z, I0_out, I2, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND0BWP7T30P140HVT (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND1BWP7T30P140HVT (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND2BWP7T30P140HVT (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX3ND4BWP7T30P140HVT (I0, I1, I2, S0, S1, ZN);
    input I0, I1, I2, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I0_out, I2, S1);
    not (ZN, I1_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D0BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D1BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D2BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4D4BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, Z);
    input I0, I1, I2, I3, S0, S1;
    output Z;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (Z, I0_out, I1_out, S1);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND0BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND1BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND2BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module MUX4ND4BWP7T30P140HVT (I0, I1, I2, I3, S0, S1, ZN);
    input I0, I1, I2, I3, S0, S1;
    output ZN;
    tsmc_mux (I0_out, I0, I1, S0);
    tsmc_mux (I1_out, I2, I3, S0);
    tsmc_mux (I2_out, I0_out, I1_out, S1);
    not (ZN, I2_out);

  specify
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b0)
    (I0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1 && S1 == 1'b0)
    (I1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b1 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I3 == 1'b0 && S0 == 1'b0 && S1 == 1'b1)
    (I2 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && S0 == 1'b1 && S1 == 1'b1)
    (I3 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b1)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S1 == 1'b0)
    (S0 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b0 && I3 == 1'b0 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b1 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b1 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b1 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b1 && I3 == 1'b0 && S0 == 1'b0)
    (S1 => ZN) = (0, 0);
    if (I0 == 1'b0 && I1 == 1'b0 && I2 == 1'b0 && I3 == 1'b1 && S0 == 1'b1)
    (S1 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D0BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D12BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D16BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D3BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2D8BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD12BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD16BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD6BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND2OPTPAD8BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    and (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D0BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D3BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D4BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3D8BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD12BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD16BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD4BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD6BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND3OPTPAD8BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    and (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D0BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D1BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D2BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D3BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D4BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ND4D8BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    and (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D0BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D12BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D16BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D3BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2D8BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD12BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD16BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD6BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR2OPTPAD8BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    or (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D0BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D3BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D4BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3D8BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD12BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD16BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD4BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD6BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR3OPTPAD8BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    or (I0_out, A1, A2, A3);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D0BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D1BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D2BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D3BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D4BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module NR4D8BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    or (I0_out, A1, A2, A3, A4);
    not (ZN, I0_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D0BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D1BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D2BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA211D4BWP7T30P140HVT (A1, A2, B, C, Z);
    input A1, A2, B, C;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B, C);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D0BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D1BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D2BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA21D4BWP7T30P140HVT (A1, A2, B, Z);
    input A1, A2, B;
    output Z;
    or (I0_out, A1, A2);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D0BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D1BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D2BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA221D4BWP7T30P140HVT (A1, A2, B1, B2, C, Z);
    input A1, A2, B1, B2, C;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out, C);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D0BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D1BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D2BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA222D4BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, Z);
    input A1, A2, B1, B2, C1, C2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (Z, I0_out, I1_out, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D0BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D1BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D2BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA22D4BWP7T30P140HVT (A1, A2, B1, B2, Z);
    input A1, A2, B1, B2;
    output Z;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D0BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D1BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D2BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA31D4BWP7T30P140HVT (A1, A2, A3, B, Z);
    input A1, A2, A3, B;
    output Z;
    or (I0_out, A1, A2, A3);
    and (Z, I0_out, B);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D0BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D1BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D2BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA32D4BWP7T30P140HVT (A1, A2, A3, B1, B2, Z);
    input A1, A2, A3, B1, B2;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D0BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D1BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D2BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OA33D4BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, Z);
    input A1, A2, A3, B1, B2, B3;
    output Z;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (Z, I0_out, I1_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D0BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D1BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D2BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211D4BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211OPTBD12BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211OPTBD1BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211OPTBD2BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211OPTBD4BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211OPTBD6BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI211OPTBD8BWP7T30P140HVT (A1, A2, B, C, ZN);
    input A1, A2, B, C;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B, C);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && C == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D0BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21D4BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21OPTBD12BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21OPTBD1BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21OPTBD2BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21OPTBD4BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21OPTBD6BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI21OPTBD8BWP7T30P140HVT (A1, A2, B, ZN);
    input A1, A2, B;
    output ZN;
    or (I0_out, A1, A2);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D0BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D1BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D2BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI221D4BWP7T30P140HVT (A1, A2, B1, B2, C, ZN);
    input A1, A2, B1, B2, C;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out, C);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0)
    (C => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1)
    (C => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D0BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D1BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D2BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI222D4BWP7T30P140HVT (A1, A2, B1, B2, C1, C2, ZN);
    input A1, A2, B1, B2, C1, C2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    or (I2_out, C1, C2);
    and (I3_out, I0_out, I1_out, I2_out);
    not (ZN, I3_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b1 && C2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0 && C2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 && C2 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 && C2 == 1'b1)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C2 == 1'b0)
    (C1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b1 && B2 == 1'b0 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0 && B2 == 1'b1 && C1 == 1'b0)
    (C2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D0BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22D4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22OPTPBD12BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22OPTPBD1BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22OPTPBD2BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22OPTPBD4BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22OPTPBD6BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI22OPTPBD8BWP7T30P140HVT (A1, A2, B1, B2, ZN);
    input A1, A2, B1, B2;
    output ZN;
    or (I0_out, A1, A2);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D0BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D1BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D2BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI31D4BWP7T30P140HVT (A1, A2, A3, B, ZN);
    input A1, A2, A3, B;
    output ZN;
    or (I0_out, A1, A2, A3);
    and (I1_out, I0_out, B);
    not (ZN, I1_out);

  specify
    (A1 => ZN) = (0, 0);
    (A2 => ZN) = (0, 0);
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (B => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (B => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (B => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D0BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D1BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D2BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI32D4BWP7T30P140HVT (A1, A2, A3, B1, B2, ZN);
    input A1, A2, A3, B1, B2;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0)
    (B2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D0BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D1BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D2BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OAI33D4BWP7T30P140HVT (A1, A2, A3, B1, B2, B3, ZN);
    input A1, A2, A3, B1, B2, B3;
    output ZN;
    or (I0_out, A1, A2, A3);
    or (I1_out, B1, B2, B3);
    and (I2_out, I0_out, I1_out);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b1 && B3 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && B1 == 1'b0 && B2 == 1'b0 && B3 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B2 == 1'b0 && B3 == 1'b0)
    (B1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B3 == 1'b0)
    (B2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1 && B1 == 1'b0 && B2 == 1'b0)
    (B3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D0BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2D8BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2OPTPAD12BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2OPTPAD1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2OPTPAD2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2OPTPAD4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR2OPTPAD8BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    or (Z, A1, A2);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D0BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D1BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D2BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D4BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR3D8BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    or (Z, A1, A2, A3);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D0BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D1BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D2BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D4BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module OR4D8BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    or (Z, A1, A2, A3, A4);

  specify
    (A1 => Z) = (0, 0);
    (A2 => Z) = (0, 0);
    (A3 => Z) = (0, 0);
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module SDFCND0BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCND4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTAD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTAD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTAD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTBD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTBD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTBD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTCD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTCD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNOPTCD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD0BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQOPTAD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQOPTAD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQOPTAD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQOPTBD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQOPTBD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCNQOPTBD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND0BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND1BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND2BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSND4BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD0BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD1BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD2BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFCSNQD4BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD0BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD1BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD2BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFD4BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND0BWP7T30P140HVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND1BWP7T30P140HVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND2BWP7T30P140HVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCND4BWP7T30P140HVT (SI, D, SE, CP, CN, Q, QN);
    input SI, D, SE, CP, CN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD0BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD1BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD2BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQD4BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQOPTBD1BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQOPTBD2BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCNQOPTBD4BWP7T30P140HVT (SI, D, SE, CP, CN, Q);
    input SI, D, SE, CP, CN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d;
        pullup (CDN);
        pullup (SDN);
        and (D1, CN_d, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        and (D1, CN, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SDFCHK, CN_D_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SDFCHK, CN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SDFCHK, CN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SDFCHK, CN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SDFCHK, nCN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SDFCHK, nCN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SDFCHK, CN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SDFCHK, CN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SDFCHK, nCN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SDFCHK, nCN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SDFCHK, nCN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SDFCHK, nCN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SDFCHK, nCN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SDFCHK, nCN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SDFCHK, CN_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SDFCHK, CN_nSE_nSI, 1'b1);
    tsmc_xbuf (CN_nD_SI_SDFCHK, CN_nD_SI, 1'b1);
    tsmc_xbuf (nCN_D_SI_SDFCHK, nCN_D_SI, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SDFCHK, nCN_nD_SI, 1'b1);
    tsmc_xbuf (CN_D_nSI_SDFCHK, CN_D_nSI, 1'b1);
    tsmc_xbuf (CN_D_SE_SDFCHK, CN_D_SE, 1'b1);
    tsmc_xbuf (CN_nD_SE_SDFCHK, CN_nD_SE, 1'b1);
    tsmc_xbuf (nCN_D_SE_SDFCHK, nCN_D_SE, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SDFCHK, nCN_nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    and (CN_D_SE_SI, CN, D, SE, SI);
    and (CN_D_nSE_SI, CN, D, nSE, SI);
    and (CN_D_nSE_nSI, CN, D, nSE, nSI);
    and (CN_nD_SE_SI, CN, nD, SE, SI);
    and (nCN_D_SE_SI, nCN, D, SE, SI);
    and (nCN_nD_SE_SI, nCN, nD, SE, SI);
    and (CN_D_SE_nSI, CN, D, SE, nSI);
    and (CN_nD_SE_nSI, CN, nD, SE, nSI);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);
    and (nCN_D_SE_nSI, nCN, D, SE, nSI);
    and (nCN_D_nSE_SI, nCN, D, nSE, SI);
    and (nCN_D_nSE_nSI, nCN, D, nSE, nSI);
    and (nCN_nD_SE_nSI, nCN, nD, SE, nSI);
    and (nCN_nD_nSE_SI, nCN, nD, nSE, SI);
    and (nCN_nD_nSE_nSI, nCN, nD, nSE, nSI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (CN_nSE_SI, CN, nSE, SI);
    and (CN_nSE_nSI, CN, nSE, nSI);
    and (CN_nD_SI, CN, nD, SI);
    and (nCN_D_SI, nCN, D, SI);
    and (nCN_nD_SI, nCN, nD, SI);
    and (CN_D_nSI, CN, D, nSI);
    and (CN_D_SE, CN, D, SE);
    and (CN_nD_SE, CN, nD, SE);
    and (nCN_D_SE, nCN, D, SE);
    and (nCN_nD_SE, nCN, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D && CN)))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND0BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND1BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND2BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSND4BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q, QN);
    input SI, D, SE, CP, CN, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD0BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD1BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD2BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKCSNQD4BWP7T30P140HVT (SI, D, SE, CP, CN, SN, Q);
    input SI, D, SE, CP, CN, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, CN_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (DS, S, D_d);
        and (D1, DS, CN_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (DS, S, D);
        and (D1, DS, CN);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CN_D_SE_SI_SN_SDFCHK, CN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_SI_nSN_SDFCHK, CN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_SN_SDFCHK, CN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_SI_nSN_SDFCHK, CN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_SN_SDFCHK, CN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSE_nSI_nSN_SDFCHK, CN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_SN_SDFCHK, CN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SI_nSN_SDFCHK, CN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_nSN_SDFCHK, CN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_nSN_SDFCHK, CN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_SN_SDFCHK, nCN_D_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SI_nSN_SDFCHK, nCN_D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_SN_SDFCHK, nCN_nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SI_nSN_SDFCHK, nCN_nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_SN_SDFCHK, CN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSI_nSN_SDFCHK, CN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_SN_SDFCHK, CN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSI_nSN_SDFCHK, CN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SN_SDFCHK, CN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SN_SDFCHK, CN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_SN_SDFCHK, nCN_D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSI_nSN_SDFCHK, nCN_D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_SN_SDFCHK, nCN_D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_SI_nSN_SDFCHK, nCN_D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_SN_SDFCHK, nCN_D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_D_nSE_nSI_nSN_SDFCHK, nCN_D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_SN_SDFCHK, nCN_nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSI_nSN_SDFCHK, nCN_nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_SN_SDFCHK, nCN_nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_SI_nSN_SDFCHK, nCN_nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_SN_SDFCHK, nCN_nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_nSE_nSI_nSN_SDFCHK, nCN_nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nSE_SI_SN_SDFCHK, CN_nSE_SI_SN, 1'b1);
    tsmc_xbuf (CN_nSE_nSI_SN_SDFCHK, CN_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (CN_nD_SI_SN_SDFCHK, CN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_SN_SDFCHK, nCN_D_SI_SN, 1'b1);
    tsmc_xbuf (nCN_D_SI_nSN_SDFCHK, nCN_D_SI_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_SN_SDFCHK, nCN_nD_SI_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SI_nSN_SDFCHK, nCN_nD_SI_nSN, 1'b1);
    tsmc_xbuf (CN_D_nSI_SN_SDFCHK, CN_D_nSI_SN, 1'b1);
    tsmc_xbuf (CN_D_nSI_nSN_SDFCHK, CN_D_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSI_nSN_SDFCHK, CN_nD_nSI_nSN, 1'b1);
    tsmc_xbuf (CN_D_SE_SN_SDFCHK, CN_D_SE_SN, 1'b1);
    tsmc_xbuf (CN_D_SE_nSN_SDFCHK, CN_D_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_nSN_SDFCHK, CN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_SE_SN_SDFCHK, CN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_SN_SDFCHK, nCN_D_SE_SN, 1'b1);
    tsmc_xbuf (nCN_D_SE_nSN_SDFCHK, nCN_D_SE_nSN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_SN_SDFCHK, nCN_nD_SE_SN, 1'b1);
    tsmc_xbuf (nCN_nD_SE_nSN_SDFCHK, nCN_nD_SE_nSN, 1'b1);
    tsmc_xbuf (CN_nD_nSE_SI_SDFCHK, CN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CN_nD_nSE_nSI_SDFCHK, CN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCN, CN);
    not (nSN, SN);
    and (CN_D_SE_SI_SN, CN, D, SE, SI, SN);
    and (CN_D_SE_SI_nSN, CN, D, SE, SI, nSN);
    and (CN_D_nSE_SI_SN, CN, D, nSE, SI, SN);
    and (CN_D_nSE_SI_nSN, CN, D, nSE, SI, nSN);
    and (CN_D_nSE_nSI_SN, CN, D, nSE, nSI, SN);
    and (CN_D_nSE_nSI_nSN, CN, D, nSE, nSI, nSN);
    and (CN_nD_SE_SI_SN, CN, nD, SE, SI, SN);
    and (CN_nD_SE_SI_nSN, CN, nD, SE, SI, nSN);
    and (CN_nD_nSE_SI_nSN, CN, nD, nSE, SI, nSN);
    and (CN_nD_nSE_nSI_nSN, CN, nD, nSE, nSI, nSN);
    and (nCN_D_SE_SI_SN, nCN, D, SE, SI, SN);
    and (nCN_D_SE_SI_nSN, nCN, D, SE, SI, nSN);
    and (nCN_nD_SE_SI_SN, nCN, nD, SE, SI, SN);
    and (nCN_nD_SE_SI_nSN, nCN, nD, SE, SI, nSN);
    and (CN_D_SE_nSI_SN, CN, D, SE, nSI, SN);
    and (CN_D_SE_nSI_nSN, CN, D, SE, nSI, nSN);
    and (CN_nD_SE_nSI_SN, CN, nD, SE, nSI, SN);
    and (CN_nD_SE_nSI_nSN, CN, nD, SE, nSI, nSN);
    and (CN_nD_nSE_SI_SN, CN, nD, nSE, SI, SN);
    and (CN_nD_nSE_nSI_SN, CN, nD, nSE, nSI, SN);
    and (nCN_D_SE_nSI_SN, nCN, D, SE, nSI, SN);
    and (nCN_D_SE_nSI_nSN, nCN, D, SE, nSI, nSN);
    and (nCN_D_nSE_SI_SN, nCN, D, nSE, SI, SN);
    and (nCN_D_nSE_SI_nSN, nCN, D, nSE, SI, nSN);
    and (nCN_D_nSE_nSI_SN, nCN, D, nSE, nSI, SN);
    and (nCN_D_nSE_nSI_nSN, nCN, D, nSE, nSI, nSN);
    and (nCN_nD_SE_nSI_SN, nCN, nD, SE, nSI, SN);
    and (nCN_nD_SE_nSI_nSN, nCN, nD, SE, nSI, nSN);
    and (nCN_nD_nSE_SI_SN, nCN, nD, nSE, SI, SN);
    and (nCN_nD_nSE_SI_nSN, nCN, nD, nSE, SI, nSN);
    and (nCN_nD_nSE_nSI_SN, nCN, nD, nSE, nSI, SN);
    and (nCN_nD_nSE_nSI_nSN, nCN, nD, nSE, nSI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (CN_nSE_SI_SN, CN, nSE, SI, SN);
    and (CN_nSE_nSI_SN, CN, nSE, nSI, SN);
    and (CN_nD_SI_SN, CN, nD, SI, SN);
    and (nCN_D_SI_SN, nCN, D, SI, SN);
    and (nCN_D_SI_nSN, nCN, D, SI, nSN);
    and (nCN_nD_SI_SN, nCN, nD, SI, SN);
    and (nCN_nD_SI_nSN, nCN, nD, SI, nSN);
    and (CN_D_nSI_SN, CN, D, nSI, SN);
    and (CN_D_nSI_nSN, CN, D, nSI, nSN);
    and (CN_nD_nSI_nSN, CN, nD, nSI, nSN);
    and (CN_D_SE_SN, CN, D, SE, SN);
    and (CN_D_SE_nSN, CN, D, SE, nSN);
    and (CN_nD_SE_nSN, CN, nD, SE, nSN);
    and (CN_nD_SE_SN, CN, nD, SE, SN);
    and (nCN_D_SE_SN, nCN, D, SE, SN);
    and (nCN_D_SE_nSN, nCN, D, SE, nSN);
    and (nCN_nD_SE_SN, nCN, nD, SE, SN);
    and (nCN_nD_SE_nSN, nCN, nD, SE, nSN);
    and (CN_nD_nSE_SI, CN, nD, nSE, SI);
    and (CN_nD_nSE_nSI, CN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, CN_d, SN_d);
      and  (SN_check, SE_int_not, CN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, CN, SN);
      and  (SN_check, SE_int_not, CN);
    `endif
    buf  (CN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (CN_DEFCHK, CN_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && CN && D) || (!(SE) && CN && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nCN_nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier,,, CP_d, CN_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_SN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, posedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, negedge CN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nCN_nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& CN_nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND0BWP7T30P140HVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND1BWP7T30P140HVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND2BWP7T30P140HVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSND4BWP7T30P140HVT (SI, D, SE, CP, SN, Q, QN);
    input SI, D, SE, CP, SN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD0BWP7T30P140HVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD1BWP7T30P140HVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD2BWP7T30P140HVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFKSNQD4BWP7T30P140HVT (SI, D, SE, CP, SN, Q);
    input SI, D, SE, CP, SN;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d, SN_d;
        pullup (CDN);
        pullup (SDN);
        not (S, SN_d);
        or (D1, S, D_d);
        tsmc_mux (D2, D1, SI_d, SE_d);
        tsmc_dff (Q_buf, D2, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        not (S, SN);
        or (D1, S, D);
        tsmc_mux (D2, D1, SI, SE);
        tsmc_dff (Q_buf, D2, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SN_SDFCHK, D_SE_SI_SN, 1'b1);
    tsmc_xbuf (D_SE_SI_nSN_SDFCHK, D_SE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_SI_SN_SDFCHK, D_nSE_SI_SN, 1'b1);
    tsmc_xbuf (D_nSE_SI_nSN_SDFCHK, D_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SN_SDFCHK, D_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSE_nSI_nSN_SDFCHK, D_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SI_SN_SDFCHK, nD_SE_SI_SN, 1'b1);
    tsmc_xbuf (nD_SE_SI_nSN_SDFCHK, nD_SE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_nSN_SDFCHK, nD_nSE_SI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_nSN_SDFCHK, nD_nSE_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_nSI_SN_SDFCHK, D_SE_nSI_SN, 1'b1);
    tsmc_xbuf (D_SE_nSI_nSN_SDFCHK, D_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SN_SDFCHK, nD_SE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SE_nSI_nSN_SDFCHK, nD_SE_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SN_SDFCHK, nD_nSE_SI_SN, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SN_SDFCHK, nD_nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nSE_SI_SN_SDFCHK, nSE_SI_SN, 1'b1);
    tsmc_xbuf (nSE_nSI_SN_SDFCHK, nSE_nSI_SN, 1'b1);
    tsmc_xbuf (nD_SI_SN_SDFCHK, nD_SI_SN, 1'b1);
    tsmc_xbuf (D_nSI_SN_SDFCHK, D_nSI_SN, 1'b1);
    tsmc_xbuf (D_nSI_nSN_SDFCHK, D_nSI_nSN, 1'b1);
    tsmc_xbuf (nD_nSI_nSN_SDFCHK, nD_nSI_nSN, 1'b1);
    tsmc_xbuf (D_SE_SN_SDFCHK, D_SE_SN, 1'b1);
    tsmc_xbuf (D_SE_nSN_SDFCHK, D_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_nSN_SDFCHK, nD_SE_nSN, 1'b1);
    tsmc_xbuf (nD_SE_SN_SDFCHK, nD_SE_SN, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nSN, SN);
    and (D_SE_SI_SN, D, SE, SI, SN);
    and (D_SE_SI_nSN, D, SE, SI, nSN);
    and (D_nSE_SI_SN, D, nSE, SI, SN);
    and (D_nSE_SI_nSN, D, nSE, SI, nSN);
    and (D_nSE_nSI_SN, D, nSE, nSI, SN);
    and (D_nSE_nSI_nSN, D, nSE, nSI, nSN);
    and (nD_SE_SI_SN, nD, SE, SI, SN);
    and (nD_SE_SI_nSN, nD, SE, SI, nSN);
    and (nD_nSE_SI_nSN, nD, nSE, SI, nSN);
    and (nD_nSE_nSI_nSN, nD, nSE, nSI, nSN);
    and (D_SE_nSI_SN, D, SE, nSI, SN);
    and (D_SE_nSI_nSN, D, SE, nSI, nSN);
    and (nD_SE_nSI_SN, nD, SE, nSI, SN);
    and (nD_SE_nSI_nSN, nD, SE, nSI, nSN);
    and (nD_nSE_SI_SN, nD, nSE, SI, SN);
    and (nD_nSE_nSI_SN, nD, nSE, nSI, SN);
    and (nSE_SI_SN, nSE, SI, SN);
    and (nSE_nSI_SN, nSE, nSI, SN);
    and (nD_SI_SN, nD, SI, SN);
    and (D_nSI_SN, D, nSI, SN);
    and (D_nSI_nSN, D, nSI, nSN);
    and (nD_nSI_nSN, nD, nSI, nSN);
    and (D_SE_SN, D, SE, SN);
    and (D_SE_nSN, D, SE, nSN);
    and (nD_SE_nSN, nD, SE, nSN);
    and (nD_SE_SN, nD, SE, SN);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (D_check, SE_int_not, SN_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (D_check, SE_int_not, SN);
    `endif
    buf  (SN_check, SE_int_not);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);
    tsmc_xbuf (SN_DEFCHK, SN_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D) || (!(SE) && !(D) && !(SN))))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_nSN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SN_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SN_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier,,, CP_d, SN_d);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier,,, CP_d, SN_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SN_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSI_nSN_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_nSN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SN_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_SI_SDFCHK, negedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SN , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_nSE_nSI_SDFCHK, negedge SN , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMD0BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMD1BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMD2BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMD4BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q, QN);
    input DA, DB, SA, SI, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMQD0BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMQD1BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMQD2BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFMQD4BWP7T30P140HVT (DA, DB, SA, SI, SE, CP, Q);
    input DA, DB, SA, SI, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire DA_d, DB_d, SA_d, SI_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB_d, DA_d, SA_d);
        tsmc_mux (D_i, D, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D, DB, DA, SA);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (DA_DB_SA_SE_SI_SDFCHK, DA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_SI_SDFCHK, DA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSE_nSI_SDFCHK, DA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SI_SDFCHK, DA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_SI_SDFCHK, DA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSE_nSI_SDFCHK, DA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SI_SDFCHK, DA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_SI_SDFCHK, DA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSE_nSI_SDFCHK, DA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SI_SDFCHK, DA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SI_SDFCHK, nDA_DB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SI_SDFCHK, nDA_DB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_SI_SDFCHK, nDA_DB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSE_nSI_SDFCHK, nDA_DB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SI_SDFCHK, nDA_nDB_SA_SE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SI_SDFCHK, nDA_nDB_nSA_SE_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_nSI_SDFCHK, DA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_nSI_SDFCHK, DA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_nSI_SDFCHK, DA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_nSI_SDFCHK, DA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_SI_SDFCHK, DA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_nSE_nSI_SDFCHK, DA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_nSI_SDFCHK, nDA_DB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_SI_SDFCHK, nDA_DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_nSE_nSI_SDFCHK, nDA_DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_nSI_SDFCHK, nDA_DB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_nSI_SDFCHK, nDA_nDB_SA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_SI_SDFCHK, nDA_nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_nSE_nSI_SDFCHK, nDA_nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_nSI_SDFCHK, nDA_nDB_nSA_SE_nSI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_SI_SDFCHK, nDA_nDB_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_nSE_nSI_SDFCHK, nDA_nDB_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_SI_SDFCHK, DB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (DB_SA_nSE_nSI_SDFCHK, DB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_SI_SDFCHK, nDB_SA_nSE_SI, 1'b1);
    tsmc_xbuf (nDB_SA_nSE_nSI_SDFCHK, nDB_SA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_SI_SDFCHK, DA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nSA_nSE_nSI_SDFCHK, DA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_SI_SDFCHK, nDA_nSA_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_nSA_nSE_nSI_SDFCHK, nDA_nSA_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_SI_SDFCHK, DA_nDB_nSE_SI, 1'b1);
    tsmc_xbuf (DA_nDB_nSE_nSI_SDFCHK, DA_nDB_nSE_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_SI_SDFCHK, nDA_DB_nSE_SI, 1'b1);
    tsmc_xbuf (nDA_DB_nSE_nSI_SDFCHK, nDA_DB_nSE_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SI_SDFCHK, DA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SI_SDFCHK, nDA_DB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SI_SDFCHK, nDA_nDB_SA_SI, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SI_SDFCHK, nDA_nDB_nSA_SI, 1'b1);
    tsmc_xbuf (DA_DB_SA_nSI_SDFCHK, DA_DB_SA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_nSA_nSI_SDFCHK, DA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_nDB_SA_nSI_SDFCHK, DA_nDB_SA_nSI, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_nSI_SDFCHK, nDA_DB_nSA_nSI, 1'b1);
    tsmc_xbuf (DA_DB_SA_SE_SDFCHK, DA_DB_SA_SE, 1'b1);
    tsmc_xbuf (DA_DB_nSA_SE_SDFCHK, DA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_SA_SE_SDFCHK, DA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_nSA_SE_SDFCHK, nDA_DB_nSA_SE, 1'b1);
    tsmc_xbuf (DA_nDB_nSA_SE_SDFCHK, DA_nDB_nSA_SE, 1'b1);
    tsmc_xbuf (nDA_DB_SA_SE_SDFCHK, nDA_DB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_SA_SE_SDFCHK, nDA_nDB_SA_SE, 1'b1);
    tsmc_xbuf (nDA_nDB_nSA_SE_SDFCHK, nDA_nDB_nSA_SE, 1'b1);
    not (nDA, DA);
    not (nDB, DB);
    not (nSA, SA);
    not (nSI, SI);
    not (nSE, SE);
    and (DA_DB_SA_SE_SI, DA, DB, SA, SE, SI);
    and (DA_DB_SA_nSE_SI, DA, DB, SA, nSE, SI);
    and (DA_DB_SA_nSE_nSI, DA, DB, SA, nSE, nSI);
    and (DA_DB_nSA_SE_SI, DA, DB, nSA, SE, SI);
    and (DA_DB_nSA_nSE_SI, DA, DB, nSA, nSE, SI);
    and (DA_DB_nSA_nSE_nSI, DA, DB, nSA, nSE, nSI);
    and (DA_nDB_SA_SE_SI, DA, nDB, SA, SE, SI);
    and (DA_nDB_SA_nSE_SI, DA, nDB, SA, nSE, SI);
    and (DA_nDB_SA_nSE_nSI, DA, nDB, SA, nSE, nSI);
    and (DA_nDB_nSA_SE_SI, DA, nDB, nSA, SE, SI);
    and (nDA_DB_SA_SE_SI, nDA, DB, SA, SE, SI);
    and (nDA_DB_nSA_SE_SI, nDA, DB, nSA, SE, SI);
    and (nDA_DB_nSA_nSE_SI, nDA, DB, nSA, nSE, SI);
    and (nDA_DB_nSA_nSE_nSI, nDA, DB, nSA, nSE, nSI);
    and (nDA_nDB_SA_SE_SI, nDA, nDB, SA, SE, SI);
    and (nDA_nDB_nSA_SE_SI, nDA, nDB, nSA, SE, SI);
    and (DA_DB_SA_SE_nSI, DA, DB, SA, SE, nSI);
    and (DA_DB_nSA_SE_nSI, DA, DB, nSA, SE, nSI);
    and (DA_nDB_SA_SE_nSI, DA, nDB, SA, SE, nSI);
    and (DA_nDB_nSA_SE_nSI, DA, nDB, nSA, SE, nSI);
    and (DA_nDB_nSA_nSE_SI, DA, nDB, nSA, nSE, SI);
    and (DA_nDB_nSA_nSE_nSI, DA, nDB, nSA, nSE, nSI);
    and (nDA_DB_SA_SE_nSI, nDA, DB, SA, SE, nSI);
    and (nDA_DB_SA_nSE_SI, nDA, DB, SA, nSE, SI);
    and (nDA_DB_SA_nSE_nSI, nDA, DB, SA, nSE, nSI);
    and (nDA_DB_nSA_SE_nSI, nDA, DB, nSA, SE, nSI);
    and (nDA_nDB_SA_SE_nSI, nDA, nDB, SA, SE, nSI);
    and (nDA_nDB_SA_nSE_SI, nDA, nDB, SA, nSE, SI);
    and (nDA_nDB_SA_nSE_nSI, nDA, nDB, SA, nSE, nSI);
    and (nDA_nDB_nSA_SE_nSI, nDA, nDB, nSA, SE, nSI);
    and (nDA_nDB_nSA_nSE_SI, nDA, nDB, nSA, nSE, SI);
    and (nDA_nDB_nSA_nSE_nSI, nDA, nDB, nSA, nSE, nSI);
    and (DB_SA_nSE_SI, DB, SA, nSE, SI);
    and (DB_SA_nSE_nSI, DB, SA, nSE, nSI);
    and (nDB_SA_nSE_SI, nDB, SA, nSE, SI);
    and (nDB_SA_nSE_nSI, nDB, SA, nSE, nSI);
    and (DA_nSA_nSE_SI, DA, nSA, nSE, SI);
    and (DA_nSA_nSE_nSI, DA, nSA, nSE, nSI);
    and (nDA_nSA_nSE_SI, nDA, nSA, nSE, SI);
    and (nDA_nSA_nSE_nSI, nDA, nSA, nSE, nSI);
    and (DA_nDB_nSE_SI, DA, nDB, nSE, SI);
    and (DA_nDB_nSE_nSI, DA, nDB, nSE, nSI);
    and (nDA_DB_nSE_SI, nDA, DB, nSE, SI);
    and (nDA_DB_nSE_nSI, nDA, DB, nSE, nSI);
    and (DA_nDB_nSA_SI, DA, nDB, nSA, SI);
    and (nDA_DB_SA_SI, nDA, DB, SA, SI);
    and (nDA_nDB_SA_SI, nDA, nDB, SA, SI);
    and (nDA_nDB_nSA_SI, nDA, nDB, nSA, SI);
    and (DA_DB_SA_nSI, DA, DB, SA, nSI);
    and (DA_DB_nSA_nSI, DA, DB, nSA, nSI);
    and (DA_nDB_SA_nSI, DA, nDB, SA, nSI);
    and (nDA_DB_nSA_nSI, nDA, DB, nSA, nSI);
    and (DA_DB_SA_SE, DA, DB, SA, SE);
    and (DA_DB_nSA_SE, DA, DB, nSA, SE);
    and (DA_nDB_SA_SE, DA, nDB, SA, SE);
    and (nDA_DB_nSA_SE, nDA, DB, nSA, SE);
    and (DA_nDB_nSA_SE, DA, nDB, nSA, SE);
    and (nDA_DB_SA_SE, nDA, DB, SA, SE);
    and (nDA_nDB_SA_SE, nDA, nDB, SA, SE);
    and (nDA_nDB_nSA_SE, nDA, nDB, nSA, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SA_int_not, SA_d);
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
      and  (DA_check, SA_d, SE_int_not);
    `else
      not  (SA_int_not, SA);
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
      and  (DA_check, SA, SE_int_not);
    `endif
    buf  (SA_check, SE_int_not);
    and  (DB_check, SA_int_not, SE_int_not);
    or   (CP_check, SI_check, DA_check, SA_check, DB_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (DB_DEFCHK, DB_check, 1'b1);
    tsmc_xbuf (DA_DEFCHK, DA_check, 1'b1);
    tsmc_xbuf (SA_DEFCHK, SA_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && SA && DA) || (!(SE) && !(SA) && DB)))) = (0, 0);
    $width (posedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& DA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_DB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_SA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nDA_nDB_nSA_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier,,, CP_d, DA_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier,,, CP_d, DB_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier,,, CP_d, SA_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_SI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, posedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDB_SA_nSE_nSI_SDFCHK, negedge DA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_SI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, posedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nSA_nSE_nSI_SDFCHK, negedge DB , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_SI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, posedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSE_nSI_SDFCHK, negedge SA , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& DA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_DB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_SA_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nDA_nDB_nSA_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND0BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND1BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND2BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCND4BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND0BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND1BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND2BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNCSND4BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND0BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND1BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND2BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFND4BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND0BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND1BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND2BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSND4BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNCND1BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNCND2BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNCND4BWP7T30P140HVT (SI, D, SE, CPN, CDN, Q, QN);
    input SI, D, SE, CPN, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CPN_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, negedge CPN &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, negedge CPN &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, negedge CPN &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, negedge CPN &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNCSND1BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNCSND2BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNCSND4BWP7T30P140HVT (SI, D, SE, CPN, CDN, SDN, Q, QN);
    input SI, D, SE, CPN, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CPN_D_SDN_SE_SI_SDFCHK, CPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_SE_nSI_SDFCHK, CPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_SI_SDFCHK, CPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SDN_nSE_nSI_SDFCHK, CPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_SI_SDFCHK, CPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_SE_nSI_SDFCHK, CPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_SI_SDFCHK, CPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_SDN_nSE_nSI_SDFCHK, CPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_SI_SDFCHK, nCPN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_SE_nSI_SDFCHK, nCPN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_SI_SDFCHK, nCPN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SDN_nSE_nSI_SDFCHK, nCPN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_SI_SDFCHK, nCPN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_SE_nSI_SDFCHK, nCPN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_SI_SDFCHK, nCPN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SDN_nSE_nSI_SDFCHK, nCPN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_SI_SDFCHK, CDN_CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_SI_SDFCHK, CDN_CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_nSE_nSI_SDFCHK, CDN_CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_SI_SDFCHK, CDN_CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_D_SE_nSI_SDFCHK, CDN_CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_SE_nSI_SDFCHK, CDN_CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_SI_SDFCHK, CDN_CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CPN_nD_nSE_nSI_SDFCHK, CDN_CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_SI_SDFCHK, CDN_nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_SE_nSI_SDFCHK, CDN_nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_SI_SDFCHK, CDN_nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_D_nSE_nSI_SDFCHK, CDN_nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_SI_SDFCHK, CDN_nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_SE_nSI_SDFCHK, CDN_nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_SI_SDFCHK, CDN_nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCPN_nD_nSE_nSI_SDFCHK, CDN_nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (CPN_D_SDN_SE_SI, CPN, D, SDN, SE, SI);
    and (CPN_D_SDN_SE_nSI, CPN, D, SDN, SE, nSI);
    and (CPN_D_SDN_nSE_SI, CPN, D, SDN, nSE, SI);
    and (CPN_D_SDN_nSE_nSI, CPN, D, SDN, nSE, nSI);
    and (CPN_nD_SDN_SE_SI, CPN, nD, SDN, SE, SI);
    and (CPN_nD_SDN_SE_nSI, CPN, nD, SDN, SE, nSI);
    and (CPN_nD_SDN_nSE_SI, CPN, nD, SDN, nSE, SI);
    and (CPN_nD_SDN_nSE_nSI, CPN, nD, SDN, nSE, nSI);
    and (nCPN_D_SDN_SE_SI, nCPN, D, SDN, SE, SI);
    and (nCPN_D_SDN_SE_nSI, nCPN, D, SDN, SE, nSI);
    and (nCPN_D_SDN_nSE_SI, nCPN, D, SDN, nSE, SI);
    and (nCPN_D_SDN_nSE_nSI, nCPN, D, SDN, nSE, nSI);
    and (nCPN_nD_SDN_SE_SI, nCPN, nD, SDN, SE, SI);
    and (nCPN_nD_SDN_SE_nSI, nCPN, nD, SDN, SE, nSI);
    and (nCPN_nD_SDN_nSE_SI, nCPN, nD, SDN, nSE, SI);
    and (nCPN_nD_SDN_nSE_nSI, nCPN, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CPN_D_SE_SI, CDN, CPN, D, SE, SI);
    and (CDN_CPN_D_nSE_SI, CDN, CPN, D, nSE, SI);
    and (CDN_CPN_D_nSE_nSI, CDN, CPN, D, nSE, nSI);
    and (CDN_CPN_nD_SE_SI, CDN, CPN, nD, SE, SI);
    and (CDN_CPN_D_SE_nSI, CDN, CPN, D, SE, nSI);
    and (CDN_CPN_nD_SE_nSI, CDN, CPN, nD, SE, nSI);
    and (CDN_CPN_nD_nSE_SI, CDN, CPN, nD, nSE, SI);
    and (CDN_CPN_nD_nSE_nSI, CDN, CPN, nD, nSE, nSI);
    and (CDN_nCPN_D_SE_SI, CDN, nCPN, D, SE, SI);
    and (CDN_nCPN_D_SE_nSI, CDN, nCPN, D, SE, nSI);
    and (CDN_nCPN_D_nSE_SI, CDN, nCPN, D, nSE, SI);
    and (CDN_nCPN_D_nSE_nSI, CDN, nCPN, D, nSE, nSI);
    and (CDN_nCPN_nD_SE_SI, CDN, nCPN, nD, SE, SI);
    and (CDN_nCPN_nD_SE_nSI, CDN, nCPN, nD, SE, nSI);
    and (CDN_nCPN_nD_nSE_SI, CDN, nCPN, nD, nSE, SI);
    and (CDN_nCPN_nD_nSE_nSI, CDN, nCPN, nD, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CPN_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCPN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCPN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, negedge CPN &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYND1BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYND2BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYND4BWP7T30P140HVT (SI, D, SE, CPN, Q, QN);
    input SI, D, SE, CPN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CPN_check);
    pullup  (SE_check);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
  `else
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNSND1BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNSND2BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFNSYNSND4BWP7T30P140HVT (SI, D, SE, CPN, SDN, Q, QN);
    input SI, D, SE, CPN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CPN_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        not (CP, CPN_d);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        not (CP, CPN);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_D_SE_SI_SDFCHK, CPN_D_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_SI_SDFCHK, CPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_D_nSE_nSI_SDFCHK, CPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_SI_SDFCHK, CPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CPN_D_SE_nSI_SDFCHK, CPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_SE_nSI_SDFCHK, CPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_SI_SDFCHK, CPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CPN_nD_nSE_nSI_SDFCHK, CPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_SI_SDFCHK, nCPN_D_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_SE_nSI_SDFCHK, nCPN_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_SI_SDFCHK, nCPN_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_D_nSE_nSI_SDFCHK, nCPN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_SI_SDFCHK, nCPN_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_SE_nSI_SDFCHK, nCPN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_SI_SDFCHK, nCPN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCPN_nD_nSE_nSI_SDFCHK, nCPN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCPN, CPN);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CPN_D_SE_SI, CPN, D, SE, SI);
    and (CPN_D_nSE_SI, CPN, D, nSE, SI);
    and (CPN_D_nSE_nSI, CPN, D, nSE, nSI);
    and (CPN_nD_SE_SI, CPN, nD, SE, SI);
    and (CPN_D_SE_nSI, CPN, D, SE, nSI);
    and (CPN_nD_SE_nSI, CPN, nD, SE, nSI);
    and (CPN_nD_nSE_SI, CPN, nD, nSE, SI);
    and (CPN_nD_nSE_nSI, CPN, nD, nSE, nSI);
    and (nCPN_D_SE_SI, nCPN, D, SE, SI);
    and (nCPN_D_SE_nSI, nCPN, D, SE, nSI);
    and (nCPN_D_nSE_SI, nCPN, D, nSE, SI);
    and (nCPN_D_nSE_nSI, nCPN, D, nSE, nSI);
    and (nCPN_nD_SE_SI, nCPN, nD, SE, SI);
    and (nCPN_nD_SE_nSI, nCPN, nD, SE, nSI);
    and (nCPN_nD_nSE_SI, nCPN, nD, nSE, SI);
    and (nCPN_nD_nSE_nSI, nCPN, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CPN_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CPN_DEFCHK, CPN_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (negedge CPN => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (negedge CPN => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CPN == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CPN &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCPN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CPN_d);
    `else
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CPN_d, D_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CPN_d, SE_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CPN_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (negedge CPN &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, negedge CPN &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, negedge CPN &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, negedge CPN &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, negedge CPN &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (negedge CPN &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (negedge CPN &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFOPTAD1BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFOPTAD2BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFOPTAD4BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFOPTBD1BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFOPTBD2BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFOPTBD4BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD0BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD1BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD2BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQD4BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND0BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND1BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND2BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQND4BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQNOPTBD1BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQNOPTBD2BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQNOPTBD4BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQOPTAD1BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQOPTAD2BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQOPTAD4BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQOPTBD1BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQOPTBD2BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFQOPTBD4BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND0BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND1BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND2BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSND4BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNOPTBD1BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNOPTBD2BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNOPTBD4BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD0BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD1BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD2BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQD4BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQOPTBD1BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQOPTBD2BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSNQOPTBD4BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCND1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCND2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCND4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q, QN);
    input SI, D, SE, CP, CDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCNQD1BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCNQD2BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCNQD4BWP7T30P140HVT (SI, D, SE, CP, CDN, Q);
    input SI, D, SE, CP, CDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d;
            buf (CDN_i, CDN_d);
        `else 
            buf (CDN_i, CDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SI_SDFCHK, CDN_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_SI_SDFCHK, CDN_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSE_nSI_SDFCHK, CDN_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SI_SDFCHK, CDN_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nSE_SI_SDFCHK, CDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nSE_nSI_SDFCHK, CDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SI_SDFCHK, CDN_nD_SI, 1'b1);
    tsmc_xbuf (CDN_D_nSI_SDFCHK, CDN_D_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SE_SDFCHK, CDN_D_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SE_SDFCHK, CDN_nD_SE, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_D_SE_SI, CDN, D, SE, SI);
    and (CDN_D_nSE_SI, CDN, D, nSE, SI);
    and (CDN_D_nSE_nSI, CDN, D, nSE, nSI);
    and (CDN_nD_SE_SI, CDN, nD, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);
    and (CDN_nSE_SI, CDN, nSE, SI);
    and (CDN_nSE_nSI, CDN, nSE, nSI);
    and (CDN_nD_SI, CDN, nD, SI);
    and (CDN_D_nSI, CDN, D, nSI);
    and (CDN_D_SE, CDN, D, SE);
    and (CDN_nD_SE, CDN, nD, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SE);
    `endif
    and  (D_check, CDN_i, SE_int_not);
    buf  (CP_check, CDN_i);
    buf  (SE_check, CDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (negedge CDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SE_SI_SDFCHK, posedge CP &&& D_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_SI_SDFCHK, posedge CP &&& D_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_nSE_nSI_SDFCHK, posedge CP &&& D_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SE_SI_SDFCHK, posedge CP &&& nD_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_SI_SDFCHK, posedge CDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCSND1BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCSND2BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCSND4BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q, QN);
    input SI, D, SE, CP, CDN, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN_buf, Q_buf);
        and (QN, QN_buf, SDN_i);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (QN-:1'b0)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (SDN => QN) = (0, 0);
    if (CDN == 1'b0 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (SDN => QN) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCSNQD1BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCSNQD2BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNCSNQD4BWP7T30P140HVT (SI, D, SE, CP, CDN, SDN, Q);
    input SI, D, SE, CP, CDN, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire CDN_d, SDN_d;
            buf (CDN_i, CDN_d);
            buf (SDN_i, SDN_d);
        `else 
            buf (CDN_i, CDN);
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (CDN_i, CDN);
        buf (SDN_i, SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN_i, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 
    `ifdef TETRAMAX
    `else
    reg flag;
    always @(CDN_i or SDN_i) begin
        if (!$test$plusargs("cdn_sdn_check_off")) begin
            flag=((CDN_i===1'b0)&&(SDN_i===1'b0));
            if (flag == 1) begin 
                if (CDN_i!==1'b0) begin
                    $display("%m > CDN is released at time %.2fns.", $realtime);
                end 
                if (SDN_i!==1'b0) begin
                    $display("%m > SDN is released at time %.2fns.", $realtime);
                end 
            end 
            if (flag == 1) begin
                $display("%m > Both CDN and SDN are enabled at time %.2fns.", $realtime);
            end 
        end 
    end 

    tsmc_xbuf (CP_D_SDN_SE_SI_SDFCHK, CP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_SE_nSI_SDFCHK, CP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_SI_SDFCHK, CP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_SDN_nSE_nSI_SDFCHK, CP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_SI_SDFCHK, CP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_SE_nSI_SDFCHK, CP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_SI_SDFCHK, CP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SDN_nSE_nSI_SDFCHK, CP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_SI_SDFCHK, nCP_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_SE_nSI_SDFCHK, nCP_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_SI_SDFCHK, nCP_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SDN_nSE_nSI_SDFCHK, nCP_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_SI_SDFCHK, nCP_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_SE_nSI_SDFCHK, nCP_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_SI_SDFCHK, nCP_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_SDN_nSE_nSI_SDFCHK, nCP_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SI_SDFCHK, CDN_D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_SI_SDFCHK, CDN_D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSE_nSI_SDFCHK, CDN_D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SI_SDFCHK, CDN_nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_nSI_SDFCHK, CDN_D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_nSI_SDFCHK, CDN_nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_SI_SDFCHK, CDN_nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_nSE_nSI_SDFCHK, CDN_nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_SI_SDFCHK, CDN_CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_SE_nSI_SDFCHK, CDN_CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_SI_SDFCHK, CDN_CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_D_nSE_nSI_SDFCHK, CDN_CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_SI_SDFCHK, CDN_CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_SE_nSI_SDFCHK, CDN_CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_SI_SDFCHK, CDN_CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_CP_nD_nSE_nSI_SDFCHK, CDN_CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_SI_SDFCHK, CDN_nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_SI_SDFCHK, CDN_nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_nSE_nSI_SDFCHK, CDN_nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_SI_SDFCHK, CDN_nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_D_SE_nSI_SDFCHK, CDN_nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_SE_nSI_SDFCHK, CDN_nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_SI_SDFCHK, CDN_nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nCP_nD_nSE_nSI_SDFCHK, CDN_nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_SI_SDFCHK, CDN_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_SDN_nSE_nSI_SDFCHK, CDN_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SI_SDFCHK, CDN_nD_SDN_SI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_nSI_SDFCHK, CDN_D_SDN_nSI, 1'b1);
    tsmc_xbuf (CDN_D_SDN_SE_SDFCHK, CDN_D_SDN_SE, 1'b1);
    tsmc_xbuf (CDN_nD_SDN_SE_SDFCHK, CDN_nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (CDN_D_SE_nSI_SDFCHK, CDN_D_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_SE_nSI_SDFCHK, CDN_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_SI_SDFCHK, CDN_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CDN_nD_nSE_nSI_SDFCHK, CDN_nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (CP_D_SDN_SE_SI, CP, D, SDN, SE, SI);
    and (CP_D_SDN_SE_nSI, CP, D, SDN, SE, nSI);
    and (CP_D_SDN_nSE_SI, CP, D, SDN, nSE, SI);
    and (CP_D_SDN_nSE_nSI, CP, D, SDN, nSE, nSI);
    and (CP_nD_SDN_SE_SI, CP, nD, SDN, SE, SI);
    and (CP_nD_SDN_SE_nSI, CP, nD, SDN, SE, nSI);
    and (CP_nD_SDN_nSE_SI, CP, nD, SDN, nSE, SI);
    and (CP_nD_SDN_nSE_nSI, CP, nD, SDN, nSE, nSI);
    and (nCP_D_SDN_SE_SI, nCP, D, SDN, SE, SI);
    and (nCP_D_SDN_SE_nSI, nCP, D, SDN, SE, nSI);
    and (nCP_D_SDN_nSE_SI, nCP, D, SDN, nSE, SI);
    and (nCP_D_SDN_nSE_nSI, nCP, D, SDN, nSE, nSI);
    and (nCP_nD_SDN_SE_SI, nCP, nD, SDN, SE, SI);
    and (nCP_nD_SDN_SE_nSI, nCP, nD, SDN, SE, nSI);
    and (nCP_nD_SDN_nSE_SI, nCP, nD, SDN, nSE, SI);
    and (nCP_nD_SDN_nSE_nSI, nCP, nD, SDN, nSE, nSI);
    and (CDN_D_SDN_SE_SI, CDN, D, SDN, SE, SI);
    and (CDN_D_SDN_nSE_SI, CDN, D, SDN, nSE, SI);
    and (CDN_D_SDN_nSE_nSI, CDN, D, SDN, nSE, nSI);
    and (CDN_nD_SDN_SE_SI, CDN, nD, SDN, SE, SI);
    and (CDN_D_SDN_SE_nSI, CDN, D, SDN, SE, nSI);
    and (CDN_nD_SDN_SE_nSI, CDN, nD, SDN, SE, nSI);
    and (CDN_nD_SDN_nSE_SI, CDN, nD, SDN, nSE, SI);
    and (CDN_nD_SDN_nSE_nSI, CDN, nD, SDN, nSE, nSI);
    and (CDN_CP_D_SE_SI, CDN, CP, D, SE, SI);
    and (CDN_CP_D_SE_nSI, CDN, CP, D, SE, nSI);
    and (CDN_CP_D_nSE_SI, CDN, CP, D, nSE, SI);
    and (CDN_CP_D_nSE_nSI, CDN, CP, D, nSE, nSI);
    and (CDN_CP_nD_SE_SI, CDN, CP, nD, SE, SI);
    and (CDN_CP_nD_SE_nSI, CDN, CP, nD, SE, nSI);
    and (CDN_CP_nD_nSE_SI, CDN, CP, nD, nSE, SI);
    and (CDN_CP_nD_nSE_nSI, CDN, CP, nD, nSE, nSI);
    and (CDN_nCP_D_SE_SI, CDN, nCP, D, SE, SI);
    and (CDN_nCP_D_nSE_SI, CDN, nCP, D, nSE, SI);
    and (CDN_nCP_D_nSE_nSI, CDN, nCP, D, nSE, nSI);
    and (CDN_nCP_nD_SE_SI, CDN, nCP, nD, SE, SI);
    and (CDN_nCP_D_SE_nSI, CDN, nCP, D, SE, nSI);
    and (CDN_nCP_nD_SE_nSI, CDN, nCP, nD, SE, nSI);
    and (CDN_nCP_nD_nSE_SI, CDN, nCP, nD, nSE, SI);
    and (CDN_nCP_nD_nSE_nSI, CDN, nCP, nD, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (CDN_SDN_nSE_SI, CDN, SDN, nSE, SI);
    and (CDN_SDN_nSE_nSI, CDN, SDN, nSE, nSI);
    and (CDN_nD_SDN_SI, CDN, nD, SDN, SI);
    and (CDN_D_SDN_nSI, CDN, D, SDN, nSI);
    and (CDN_D_SDN_SE, CDN, D, SDN, SE);
    and (CDN_nD_SDN_SE, CDN, nD, SDN, SE);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (CDN_D_SE_nSI, CDN, D, SE, nSI);
    and (CDN_nD_SE_nSI, CDN, nD, SE, nSI);
    and (CDN_nD_nSE_SI, CDN, nD, nSE, SI);
    and (CDN_nD_nSE_nSI, CDN, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, CDN_i, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, CDN_i, SDN_i, SE);
    `endif
    and  (D_check, CDN_i, SDN_i, SE_int_not);
    and  (CP_check, CDN_i, SDN_i);
    and  (SE_check, CDN_i, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge CDN => (Q+:1'b0)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (CDN => Q) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SDN == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (CDN => Q) = (0, 0);
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CDN == 1'b1 && CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (negedge CDN &&& CP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& CP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CDN &&& nCP_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& CDN_nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CDN_nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0,0, notifier, , , CDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier,,, SDN_d, CDN_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier,,, CDN_d, SDN_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
      $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
      $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge SDN &&& CP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& CP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_D_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_SE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_SI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge CDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& CP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_D_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_SE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_SI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CDN &&& nCP_nD_nSE_nSI_SDFCHK, posedge SDN , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& CDN_nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_SE_SI_SDFCHK, posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_SI_SDFCHK, posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& D_SDN_nSE_nSI_SDFCHK, posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge CDN &&& nD_SDN_SE_SI_SDFCHK, posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_SI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, posedge CDN , 0, notifier);
    $hold (posedge CP &&& nD_SDN_SE_SI_SDFCHK, posedge CDN , 0, notifier);
    $recovery (posedge SDN &&& CDN_D_SE_nSI_SDFCHK, posedge CP &&& CDN_D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_SE_nSI_SDFCHK, posedge CP &&& CDN_nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_SI_SDFCHK, posedge CP &&& CDN_nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& CDN_nD_nSE_nSI_SDFCHK, posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& CDN_D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& CDN_nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYND1BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYND2BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYND4BWP7T30P140HVT (SI, D, SE, CP, Q, QN);
    input SI, D, SE, CP;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNQD1BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNQD2BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNQD4BWP7T30P140HVT (SI, D, SE, CP, Q);
    input SI, D, SE, CP;
    output Q;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (nD_SI, nD, SI);
    and (D_nSI, D, nSI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNQND1BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNQND2BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNQND4BWP7T30P140HVT (SI, D, SE, CP, QN);
    input SI, D, SE, CP;
    output QN;
    reg notifier;
    `ifdef NTC
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN, notifier);
        not (QN, Q_buf);
    `else 
        pullup (CDN);
        pullup (SDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN, notifier);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    tsmc_xbuf (D_SE_SI_SDFCHK, D_SE_SI, 1'b1);
    tsmc_xbuf (D_nSE_SI_SDFCHK, D_nSE_SI, 1'b1);
    tsmc_xbuf (D_nSE_nSI_SDFCHK, D_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_SI_SDFCHK, nD_SE_SI, 1'b1);
    tsmc_xbuf (nSE_SI_SDFCHK, nSE_SI, 1'b1);
    tsmc_xbuf (nSE_nSI_SDFCHK, nSE_nSI, 1'b1);
    tsmc_xbuf (D_nSI_SDFCHK, D_nSI, 1'b1);
    tsmc_xbuf (nD_SI_SDFCHK, nD_SI, 1'b1);
    tsmc_xbuf (D_SE_SDFCHK, D_SE, 1'b1);
    tsmc_xbuf (nD_SE_SDFCHK, nD_SE, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);
    and (D_SE_SI, D, SE, SI);
    and (D_nSE_SI, D, nSE, SI);
    and (D_nSE_nSI, D, nSE, nSI);
    and (nD_SE_SI, nD, SE, SI);
    and (nSE_SI, nSE, SI);
    and (nSE_nSI, nSE, nSI);
    and (D_nSI, D, nSI);
    and (nD_SI, nD, SI);
    and (D_SE, D, SE);
    and (nD_SE, nD, SE);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      buf  (SI_check, SE_d);
    `else
      not  (SE_int_not, SE);
      buf  (SI_check, SE);
    `endif
    buf  (D_check, SE_int_not);
    pullup  (CP_check);
    pullup  (SE_check);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    $width (posedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SE_SI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
  `else
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SE_SDFCHK, negedge SI , 0, 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNSND1BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNSND2BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNSND4BWP7T30P140HVT (SI, D, SE, CP, SDN, Q, QN);
    input SI, D, SE, CP, SDN;
    output Q, QN;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
        not (QN, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    (posedge CP => (QN-:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (QN-:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNSNQD1BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNSNQD2BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module SDFSYNSNQD4BWP7T30P140HVT (SI, D, SE, CP, SDN, Q);
    input SI, D, SE, CP, SDN;
    output Q;
    reg notifier;
    `ifdef NTC
        `ifdef RECREM
            wire SDN_d;
            buf (SDN_i, SDN_d);
        `else 
            buf (SDN_i, SDN);
        `endif 
        wire SI_d, D_d, SE_d, CP_d;
        pullup (CDN);
        tsmc_mux (D_i, D_d, SI_d, SE_d);
        tsmc_dff (Q_buf, D_i, CP_d, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `else 
        buf (SDN_i, SDN);
        pullup (CDN);
        tsmc_mux (D_i, D, SI, SE);
        tsmc_dff (Q_buf, D_i, CP, CDN, SDN_i, notifier);
        buf (Q, Q_buf);
    `endif 

  `ifdef TETRAMAX
  `else
    tsmc_xbuf (D_SDN_SE_SI_SDFCHK, D_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_SI_SDFCHK, D_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSE_nSI_SDFCHK, D_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SI_SDFCHK, nD_SDN_SE_SI, 1'b1);
    tsmc_xbuf (D_SDN_SE_nSI_SDFCHK, D_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SE_nSI_SDFCHK, nD_SDN_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_SI_SDFCHK, nD_SDN_nSE_SI, 1'b1);
    tsmc_xbuf (nD_SDN_nSE_nSI_SDFCHK, nD_SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_D_SE_SI_SDFCHK, CP_D_SE_SI, 1'b1);
    tsmc_xbuf (CP_D_SE_nSI_SDFCHK, CP_D_SE_nSI, 1'b1);
    tsmc_xbuf (CP_D_nSE_SI_SDFCHK, CP_D_nSE_SI, 1'b1);
    tsmc_xbuf (CP_D_nSE_nSI_SDFCHK, CP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_SE_SI_SDFCHK, CP_nD_SE_SI, 1'b1);
    tsmc_xbuf (CP_nD_SE_nSI_SDFCHK, CP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_SI_SDFCHK, CP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (CP_nD_nSE_nSI_SDFCHK, CP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_D_SE_SI_SDFCHK, nCP_D_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_SI_SDFCHK, nCP_D_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_D_nSE_nSI_SDFCHK, nCP_D_nSE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_SI_SDFCHK, nCP_nD_SE_SI, 1'b1);
    tsmc_xbuf (nCP_D_SE_nSI_SDFCHK, nCP_D_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_SE_nSI_SDFCHK, nCP_nD_SE_nSI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_SI_SDFCHK, nCP_nD_nSE_SI, 1'b1);
    tsmc_xbuf (nCP_nD_nSE_nSI_SDFCHK, nCP_nD_nSE_nSI, 1'b1);
    tsmc_xbuf (SDN_nSE_SI_SDFCHK, SDN_nSE_SI, 1'b1);
    tsmc_xbuf (SDN_nSE_nSI_SDFCHK, SDN_nSE_nSI, 1'b1);
    tsmc_xbuf (nD_SDN_SI_SDFCHK, nD_SDN_SI, 1'b1);
    tsmc_xbuf (D_SDN_nSI_SDFCHK, D_SDN_nSI, 1'b1);
    tsmc_xbuf (D_SDN_SE_SDFCHK, D_SDN_SE, 1'b1);
    tsmc_xbuf (nD_SDN_SE_SDFCHK, nD_SDN_SE, 1'b1);
    tsmc_xbuf (D_SE_nSI_SDFCHK, D_SE_nSI, 1'b1);
    tsmc_xbuf (nD_SE_nSI_SDFCHK, nD_SE_nSI, 1'b1);
    tsmc_xbuf (nD_nSE_SI_SDFCHK, nD_nSE_SI, 1'b1);
    tsmc_xbuf (nD_nSE_nSI_SDFCHK, nD_nSE_nSI, 1'b1);
    not (nSI, SI);
    not (nD, D);
    not (nSE, SE);
    not (nCP, CP);
    and (D_SDN_SE_SI, D, SDN, SE, SI);
    and (D_SDN_nSE_SI, D, SDN, nSE, SI);
    and (D_SDN_nSE_nSI, D, SDN, nSE, nSI);
    and (nD_SDN_SE_SI, nD, SDN, SE, SI);
    and (D_SDN_SE_nSI, D, SDN, SE, nSI);
    and (nD_SDN_SE_nSI, nD, SDN, SE, nSI);
    and (nD_SDN_nSE_SI, nD, SDN, nSE, SI);
    and (nD_SDN_nSE_nSI, nD, SDN, nSE, nSI);
    and (CP_D_SE_SI, CP, D, SE, SI);
    and (CP_D_SE_nSI, CP, D, SE, nSI);
    and (CP_D_nSE_SI, CP, D, nSE, SI);
    and (CP_D_nSE_nSI, CP, D, nSE, nSI);
    and (CP_nD_SE_SI, CP, nD, SE, SI);
    and (CP_nD_SE_nSI, CP, nD, SE, nSI);
    and (CP_nD_nSE_SI, CP, nD, nSE, SI);
    and (CP_nD_nSE_nSI, CP, nD, nSE, nSI);
    and (nCP_D_SE_SI, nCP, D, SE, SI);
    and (nCP_D_nSE_SI, nCP, D, nSE, SI);
    and (nCP_D_nSE_nSI, nCP, D, nSE, nSI);
    and (nCP_nD_SE_SI, nCP, nD, SE, SI);
    and (nCP_D_SE_nSI, nCP, D, SE, nSI);
    and (nCP_nD_SE_nSI, nCP, nD, SE, nSI);
    and (nCP_nD_nSE_SI, nCP, nD, nSE, SI);
    and (nCP_nD_nSE_nSI, nCP, nD, nSE, nSI);
    and (SDN_nSE_SI, SDN, nSE, SI);
    and (SDN_nSE_nSI, SDN, nSE, nSI);
    and (nD_SDN_SI, nD, SDN, SI);
    and (D_SDN_nSI, D, SDN, nSI);
    and (D_SDN_SE, D, SDN, SE);
    and (nD_SDN_SE, nD, SDN, SE);
    and (D_SE_nSI, D, SE, nSI);
    and (nD_SE_nSI, nD, SE, nSI);
    and (nD_nSE_SI, nD, nSE, SI);
    and (nD_nSE_nSI, nD, nSE, nSI);


  // Timing logics defined for default constraint check
    `ifdef NTC
      not  (SE_int_not, SE_d);
      and  (SI_check, SDN_i, SE_d);
    `else
      not  (SE_int_not, SE);
      and  (SI_check, SDN_i, SE);
    `endif
    and  (D_check, SDN_i, SE_int_not);
    buf  (CP_check, SDN_i);
    buf  (SE_check, SDN_i);
    tsmc_xbuf (CP_DEFCHK, CP_check, 1'b1);
    tsmc_xbuf (SE_DEFCHK, SE_check, 1'b1);
    tsmc_xbuf (D_DEFCHK, D_check, 1'b1);
    tsmc_xbuf (SI_DEFCHK, SI_check, 1'b1);

  specify
    (posedge CP => (Q+:((SE && SI) || (!(SE) && D)))) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b1 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b1 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b1 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b1)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    if (CP == 1'b0 && D == 1'b0 && SE == 1'b0 && SI == 1'b0)
    (negedge SDN => (Q+:1'b1)) = (0, 0);
    $width (posedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& D_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (posedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge CP &&& nD_SDN_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& CP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_nSE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_D_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_SE_nSI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_SI_SDFCHK, 0, 0, notifier);
    $width (negedge SDN &&& nCP_nD_nSE_nSI_SDFCHK, 0, 0, notifier);
  `ifdef NTC
    `ifdef RECREM
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recrem (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
      $recrem (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0,0, notifier, , , SDN_d, CP_d);
    `else
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier,,, CP_d, D_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier,,, CP_d, SE_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier,,, CP_d, SI_d);
      $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
      $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
      $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
      $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
    `endif
  `else
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_SI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, posedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& SDN_nSE_nSI_SDFCHK, negedge D , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, posedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_nSI_SDFCHK, negedge SE , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& D_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, posedge SI , 0, 0, notifier);
    $setuphold (posedge CP &&& nD_SDN_SE_SDFCHK, negedge SI , 0, 0, notifier);
    $recovery (posedge SDN &&& D_SE_nSI_SDFCHK, posedge CP &&& D_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_SE_nSI_SDFCHK, posedge CP &&& nD_SE_nSI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_SI_SDFCHK, posedge CP &&& nD_nSE_SI_SDFCHK, 0, notifier);
    $recovery (posedge SDN &&& nD_nSE_nSI_SDFCHK, posedge CP &&& nD_nSE_nSI_SDFCHK, 0, notifier);
    $hold (posedge CP &&& D_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_SE_nSI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_SI_SDFCHK, posedge SDN , 0, notifier);
    $hold (posedge CP &&& nD_nSE_nSI_SDFCHK, posedge SDN , 0, notifier);
  `endif
  endspecify
  `endif
endmodule
`endcelldefine

`celldefine
module TAPCELLBWP7T30P140;
    // No function
endmodule
`endcelldefine

`celldefine
module TIEHBWP7T30P140HVT (Z);
    output Z;
    buf (Z, 1'b1);

endmodule
`endcelldefine

`celldefine
module TIELBWP7T30P140HVT (ZN);
    output ZN;
    buf (ZN, 1'b0);

endmodule
`endcelldefine

`celldefine
module XNR2D0BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2D4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2OPTND1BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2OPTND2BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2OPTND4BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR2OPTND6BWP7T30P140HVT (A1, A2, ZN);
    input A1, A2;
    output ZN;
    xor (I0_out, A1, A2);
    not (ZN, I0_out);

  specify
    if (A2 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0)
    (A2 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D0BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3D4BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3OPTND1BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3OPTND2BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR3OPTND4BWP7T30P140HVT (A1, A2, A3, ZN);
    input A1, A2, A3;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    not (ZN, I1_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D0BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D1BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D2BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XNR4D4BWP7T30P140HVT (A1, A2, A3, A4, ZN);
    input A1, A2, A3, A4;
    output ZN;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (I2_out, I1_out, A4);
    not (ZN, I2_out);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => ZN) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => ZN) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D0BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2D4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2OPTND1BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2OPTND2BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2OPTND4BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR2OPTND6BWP7T30P140HVT (A1, A2, Z);
    input A1, A2;
    output Z;
    xor (Z, A1, A2);

  specify
    if (A2 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1)
    (A2 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D0BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D1BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D2BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3D4BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3OPTND1BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3OPTND2BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR3OPTND4BWP7T30P140HVT (A1, A2, A3, Z);
    input A1, A2, A3;
    output Z;
    xor (I0_out, A1, A2);
    xor (Z, I0_out, A3);

  specify
    if (A2 == 1'b1 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1)
    (A3 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D0BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D1BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D2BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module XOR4D4BWP7T30P140HVT (A1, A2, A3, A4, Z);
    input A1, A2, A3, A4;
    output Z;
    xor (I0_out, A1, A2);
    xor (I1_out, I0_out, A3);
    xor (Z, I1_out, A4);

  specify
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A1 => Z) = (0, 0);
    if (A2 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A1 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b1 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A3 == 1'b0 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b1 && A4 == 1'b0)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b0 && A3 == 1'b0 && A4 == 1'b1)
    (A2 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A4 == 1'b1)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A4 == 1'b0)
    (A3 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b1 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b0 && A3 == 1'b1)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b1 && A2 == 1'b0 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
    if (A1 == 1'b0 && A2 == 1'b1 && A3 == 1'b0)
    (A4 => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID1BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID2BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID4BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOHID8BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD1BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD2BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD4BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOLOD8BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOSRHID2BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOSRHID4BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOSRHID8BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    or (Z, I, ISO);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOSRLOD2BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOSRLOD4BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module ISOSRLOD8BWP7T30P140HVT (ISO, I, Z);
    input ISO, I;
    output Z;
    not (ISO1, ISO);
    nand (Z1, ISO1, I);
    not (Z, Z1);

  specify
    (I => Z) = (0, 0);
    (ISO => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCD1BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (IN, I);
    nand (Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCD2BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (IN, I);
    nand (Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCD4BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (IN, I);
    nand (Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCD8BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (IN, I);
    nand (Z, IN, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCLOD1BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCLOD2BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCLOD4BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLCLOD8BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLHLD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD1BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD2BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD4BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCD8BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCLOD1BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCLOD2BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCLOD4BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHCLOD8BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    and (Z, I, NSLEEP);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD1BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLLHD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLSRLHCD2BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLSRLHCD4BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLSRLHCD8BWP7T30P140HVT (I, NSLEEP, Z);
    input I, NSLEEP;
    output Z;
    not (NSLEEPN, NSLEEP);
    or (Z, I, NSLEEPN);

  specify
    (I => Z) = (0, 0);
    (NSLEEP => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLSRLHD2BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLSRLHD4BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

`celldefine
module LVLSRLHD8BWP7T30P140HVT (I, Z);
    input I;
    output Z;
    buf (Z, I);

  specify
    (I => Z) = (0, 0);
  endspecify
endmodule
`endcelldefine

primitive tsmc_dff (q, d, cp, cdn, sdn, notifier);
   output q;
   input d, cp, cdn, sdn, notifier;
   reg q;
   table
      ?   ?   0   ?   ? : ? : 0 ; // CDN dominate SDN
      ?   ?   1   0   ? : ? : 1 ; // SDN is set   
      ?   ?   1   x   ? : 0 : x ; // SDN affect Q
      ?   ?   1   x   ? : 1 : 1 ; // Q=1,preset=X
      ?   ?   x   1   ? : 0 : 0 ; // Q=0,clear=X
      0 (01)  ?   1   ? : ? : 0 ; // Latch 0
      0 (0x)  1   1   ? : ? : x ; // Weak clock
      0   0   ?   1   ? : 0 : 0 ; // Keep 0 (D==Q)
      1 (01)  1   ?   ? : ? : 1 ; // Latch 1   
      1 (0x)  1   ?   ? : ? : x ; // Weak clock
      1   0   1   ?   ? : 1 : 1 ; // Keep 1 (D==Q)
      ? (1?)  1   1   ? : ? : - ; // ignore negative edge of clock
      ?   0   1   1   ? : ? : - ; // ignore low-level clock
      ?   ? (?1)  1   ? : ? : - ; // ignore positive edge of CDN
      ?   ?   1 (?1)  ? : ? : - ; // ignore posative edge of SDN
      *   ?   1   1   ? : ? : - ; // ignore data change on steady clock
      ?   ?   ?   ?   * : ? : x ; // timing check violation
   endtable
endprimitive

primitive tsmc_dla (q, d, e, cdn, sdn, notifier);
   output q;
   reg q;
   input d, e, cdn, sdn, notifier;
   table
   1  1   1   ?   ?   : ?  :  1  ; // Latch 1
   0  1   ?   1   ?   : ?  :  0  ; // Latch 0
   0 (10) 1   1   ?   : ?  :  0  ; // Latch 0 after falling edge
   1 (10) 1   1   ?   : ?  :  1  ; // Latch 1 after falling edge
   *  0   ?   ?   ?   : ?  :  -  ; // no changes
   ?  ?   ?   0   ?   : ?  :  1  ; // preset to 1
   ?  0   1   *   ?   : 1  :  1  ;
   1  ?   1   *   ?   : 1  :  1  ;
   1  *   1   ?   ?   : 1  :  1  ;
   ?  ?   0   1   ?   : ?  :  0  ; // reset to 0
   ?  0   *   1   ?   : 0  :  0  ;
   0  ?   *   1   ?   : 0  :  0  ;
   0  *   ?   1   ?   : 0  :  0  ;
   ?  ?   ?   ?   *   : ?  :  x  ; // toggle notifier
   endtable
endprimitive

primitive tsmc_mux (q, d0, d1, s);
   output q;
   input s, d0, d1;

   table
   // d0  d1  s   : q 
      0   ?   0   : 0 ;
      1   ?   0   : 1 ;
      ?   0   1   : 0 ;
      ?   1   1   : 1 ;
      0   0   x   : 0 ;
      1   1   x   : 1 ;
   endtable
endprimitive

primitive tsmc_xbuf (o, i, dummy);
   output o;     
   input i, dummy;
   table         
   // i dummy : o
      0   1   : 0 ;
      1   1   : 1 ;
      x   1   : 1 ;
   endtable      
endprimitive 

